netcdf sp041_20191205T1757 {
dimensions:
	N_PARAM = 5 ;
	N_MEASUREMENTS = 25 ;
variables:
	string TRAJECTORY ;
		TRAJECTORY:cf_role = "trajectory_id" ;
		TRAJECTORY:long_name = "trajectory name" ;
		TRAJECTORY:data_mode_vocabulary = "http://vocab.nerc.ac.uk/collection/OGXXX/" ;
	string PARAMETER(N_PARAM) ;
		PARAMETER:long_name = "name of parameter computed from glider measurements" ;
		PARAMETER:parameter_vocabulary = "https://vocab.nerc.ac.uk/collection/OG1/current/" ;
		PARAMETER:coordinates = "TRAJECTORY" ;
	double TIME_GPS(N_MEASUREMENTS) ;
		TIME_GPS:_FillValue = -1. ;
		TIME_GPS:long_name = "time of each GPS location" ;
		TIME_GPS:units = "seconds since 1970-01-01T00:00:00Z" ;
		TIME_GPS:ancillary_variables = "TIME_GPS_QC" ;
		TIME_GPS:coordinates = "TRAJECTORY" ;
	byte TIME_GPS_QC(N_MEASUREMENTS) ;
		TIME_GPS_QC:_FillValue = 0b ;
		TIME_GPS_QC:long_name = "quality flag" ;
		TIME_GPS_QC:coordinates = "TRAJECTORY" ;
	double LATITUDE_GPS(N_MEASUREMENTS) ;
		LATITUDE_GPS:_FillValue = NaN ;
		LATITUDE_GPS:long_name = "latitude of each GPS location" ;
		LATITUDE_GPS:standard_name = "latitude" ;
		LATITUDE_GPS:units = "degrees_north" ;
		LATITUDE_GPS:ancillary_variables = "LATITUDE_GPS_QC" ;
		LATITUDE_GPS:valid_max = "90" ;
		LATITUDE_GPS:valid_min = "-90" ;
		LATITUDE_GPS:coordinates = "TRAJECTORY" ;
	byte LATITUDE_GPS_QC(N_MEASUREMENTS) ;
		LATITUDE_GPS_QC:_FillValue = 0b ;
		LATITUDE_GPS_QC:long_name = "quality flag" ;
		LATITUDE_GPS_QC:coordinates = "TRAJECTORY" ;
	double LONGITUDE_GPS(N_MEASUREMENTS) ;
		LONGITUDE_GPS:_FillValue = NaN ;
		LONGITUDE_GPS:long_name = "longitude of each GPS location" ;
		LONGITUDE_GPS:standard_name = "longitude" ;
		LONGITUDE_GPS:units = "degrees_east" ;
		LONGITUDE_GPS:ancillary_variables = "LONGITUDE_GPS_QC" ;
		LONGITUDE_GPS:valid_max = "180" ;
		LONGITUDE_GPS:valid_min = "-180" ;
		LONGITUDE_GPS:coordinates = "TRAJECTORY" ;
	byte LONGITUDE_GPS_QC(N_MEASUREMENTS) ;
		LONGITUDE_GPS_QC:_FillValue = 0b ;
		LONGITUDE_GPS_QC:long_name = "quality flag" ;
		LONGITUDE_GPS_QC:coordinates = "TRAJECTORY" ;
	string PLATFORM ;
		PLATFORM:coordinates = "TRAJECTORY" ;
	byte PHASE(N_MEASUREMENTS) ;
		PHASE:_FillValue = 0b ;
		PHASE:long_name = "behavior of the glider at sea" ;
		PHASE:ancillary_variables = "PHASE_QC" ;
		PHASE:phase_vocabulary = "url to phase vocab list" ;
		PHASE:phase_calculation_method = "TBD" ;
		PHASE:phase_calculation_method_vocabulary = "TBD" ;
		PHASE:phase_calculation_method_doi = "TBD" ;
		PHASE:coordinates = "TRAJECTORY" ;
	byte PHASE_QC(N_MEASUREMENTS) ;
		PHASE_QC:_FillValue = 0b ;
		PHASE_QC:long_name = "quality flag" ;
		PHASE_QC:coordinates = "TRAJECTORY" ;
	double TIME(N_MEASUREMENTS) ;
		TIME:_FillValue = -1. ;
		TIME:long_name = "time of measurement and GPS location" ;
		TIME:standard_name = "time" ;
		TIME:calendar = "gregorian" ;
		TIME:units = "seconds since 1970-01-01T00:00:00Z" ;
		TIME:coordinates = "TRAJECTORY" ;
	double LATITUDE(N_MEASUREMENTS) ;
		LATITUDE:_FillValue = -9999.9 ;
		LATITUDE:long_name = "latitude of each measurement and GPS location" ;
		LATITUDE:standard_name = "latitude" ;
		LATITUDE:units = "degrees_north" ;
		LATITUDE:valid_max = "90" ;
		LATITUDE:valid_min = "-90" ;
		LATITUDE:coordinates = "TRAJECTORY" ;
	double LONGITUDE(N_MEASUREMENTS) ;
		LONGITUDE:_FillValue = -9999.9 ;
		LONGITUDE:long_name = "longitude of each measurement and GPS location" ;
		LONGITUDE:standard_name = "longitude" ;
		LONGITUDE:units = "degrees_east" ;
		LONGITUDE:valid_max = "180" ;
		LONGITUDE:valid_min = "-180" ;
		LONGITUDE:coordinates = "TRAJECTORY" ;
	double PRES(N_MEASUREMENTS) ;
		PRES:_FillValue = -9999.9 ;
		PRES:long_name = "Pressure" ;
		PRES:standard_name = "sea_water_pressure" ;
		PRES:units = "dbar" ;
		PRES:ancillary_variables = "PRES_QC" ;
		PRES:comment = "Sea water pressure, equals 0 at sea-level" ;
		PRES:sensor = "/CTD" ;
		PRES:coordinates = "TRAJECTORY" ;
	byte PRES_QC(N_MEASUREMENTS) ;
		PRES_QC:_FillValue = 0b ;
		PRES_QC:long_name = "quality flag" ;
		PRES_QC:coordinates = "TRAJECTORY" ;
	double DEPTH(N_MEASUREMENTS) ;
		DEPTH:_FillValue = NaN ;
		DEPTH:long_name = "Depth" ;
		DEPTH:standard_name = "depth" ;
		DEPTH:units = "m" ;
		DEPTH:positive = "down" ;
		DEPTH:sensor = "/CTD" ;
		DEPTH:coordinates = "TRAJECTORY" ;
	double TEMP(N_MEASUREMENTS) ;
		TEMP:_FillValue = -9999.9 ;
		TEMP:long_name = "Sea Water Temperature" ;
		TEMP:standard_name = "sea_water_temperature" ;
		TEMP:units = "Celsius" ;
		TEMP:ancillary_variables = "TEMP_QC" ;
		TEMP:valid_max = 40. ;
		TEMP:valid_min = -5. ;
		TEMP:coverage_content_type = "physicalMeasurement" ;
		TEMP:coordinates = "time lon lat depth" ;
		TEMP:comment = "Sea temperature in-situ ITS-90 scale" ;
		TEMP:sensor = "/CTD" ;
	byte TEMP_QC(N_MEASUREMENTS) ;
		TEMP_QC:_FillValue = 0b ;
		TEMP_QC:long_name = "quality flag" ;
		TEMP_QC:coordinates = "TRAJECTORY" ;
	double PSAL(N_MEASUREMENTS) ;
		PSAL:_FillValue = NaN ;
		PSAL:long_name = "Sea Water Salinity" ;
		PSAL:standard_name = "sea_water_practical_salinity" ;
		PSAL:units = "1" ;
		PSAL:ancillary_variables = "PSAL_QC" ;
		PSAL:valid_max = 40. ;
		PSAL:valid_min = 0. ;
		PSAL:coverage_content_type = "physicalMeasurement" ;
		PSAL:coordinates = "time lon lat depth" ;
		PSAL:comment = "Practical salinity computed using UNESCO 1983 algorithm" ;
		PSAL:sensor = "/CTD" ;
	byte PSAL_QC(N_MEASUREMENTS) ;
		PSAL_QC:_FillValue = 0b ;
		PSAL_QC:long_name = "quality flag" ;
		PSAL_QC:coordinates = "TRAJECTORY" ;
	double DEPLOYMENT_TIME ;
		DEPLOYMENT_TIME:_FillValue = -1. ;
		DEPLOYMENT_TIME:long_name = "date of deployment" ;
		DEPLOYMENT_TIME:standard_name = "time" ;
		DEPLOYMENT_TIME:calendar = "gregorian" ;
		DEPLOYMENT_TIME:units = "seconds since 1970-01-01T00:00:00Z" ;
		DEPLOYMENT_TIME:coordinates = "TRAJECTORY" ;
	double DEPLOYMENT_LATITUDE ;
		DEPLOYMENT_LATITUDE:_FillValue = NaN ;
		DEPLOYMENT_LATITUDE:long_name = "latitude of deployment" ;
		DEPLOYMENT_LATITUDE:standard_name = "latitude" ;
		DEPLOYMENT_LATITUDE:units = "degrees_north" ;
		DEPLOYMENT_LATITUDE:valid_max = "90" ;
		DEPLOYMENT_LATITUDE:valid_min = "-90" ;
		DEPLOYMENT_LATITUDE:coordinates = "TRAJECTORY" ;
	double DEPLOYMENT_LONGITUDE ;
		DEPLOYMENT_LONGITUDE:_FillValue = NaN ;
		DEPLOYMENT_LONGITUDE:long_name = "longitude of deployment" ;
		DEPLOYMENT_LONGITUDE:standard_name = "longitude" ;
		DEPLOYMENT_LONGITUDE:units = "degrees_east" ;
		DEPLOYMENT_LONGITUDE:valid_max = "180" ;
		DEPLOYMENT_LONGITUDE:valid_min = "-180" ;
		DEPLOYMENT_LONGITUDE:coordinates = "TRAJECTORY" ;
	string TELECOM_TYPE ;
		TELECOM_TYPE:long_name = "type of telecommunication systems used by the glider" ;
		TELECOM_TYPE:telecom_type_vocabulary = "TBD" ;
		TELECOM_TYPE:coordinates = "TRAJECTORY" ;
	string TRACKING_SYSTEM ;
		TRACKING_SYSTEM:long_name = "type of tracking systems used by the glider" ;
		TRACKING_SYSTEM:tracking_system_vocabulary = "TBD" ;
		TRACKING_SYSTEM:coordinates = "TRAJECTORY" ;
	int N_MEASUREMENTS(N_MEASUREMENTS) ;
	string PLATFORM_TYPE ;
		PLATFORM_TYPE:long_name = "type of glider" ;
		PLATFORM_TYPE:platform_type_vocabulary = "https://vocab.nerc.ac.uk/collection/L06/current/" ;
		PLATFORM_TYPE:coordinates = "TRAJECTORY" ;
	string PLATFORM_MODEL ;
		PLATFORM_MODEL:long_name = "model of the glider" ;
		PLATFORM_MODEL:platform_model_vocabulary = "http://vocab.nerc.ac.uk/collection/B76/current/B7600027/" ;
		PLATFORM_MODEL:coordinates = "TRAJECTORY" ;
	string PLATFORM_MAKER ;
		PLATFORM_MAKER:long_name = "Glider manufacturer" ;
		PLATFORM_MAKER:platform_maker_vocabulary = "TBD" ;
		PLATFORM_MAKER:coordinates = "TRAJECTORY" ;
	string PLATFORM_SERIAL_NUMBER ;
		PLATFORM_SERIAL_NUMBER:long_name = "glider serial number" ;
		PLATFORM_SERIAL_NUMBER:coordinates = "TRAJECTORY" ;
	string PLATFORM_CODE ;
		PLATFORM_CODE:long_name = "nickname of the glider" ;
		PLATFORM_CODE:coordinates = "TRAJECTORY" ;
	int PLATFORM_DEPTH_RATING ;
		PLATFORM_DEPTH_RATING:long_name = "Depth limit in meters of the glider for this mission" ;
		PLATFORM_DEPTH_RATING:coordinates = "TRAJECTORY" ;
	string WMO_IDENTIFIER ;
		WMO_IDENTIFIER:long_name = "wmo id" ;
		WMO_IDENTIFIER:coordinates = "TRAJECTORY" ;

// global attributes:
		:Conventions = "CF-1.8, ACDD-1.3, OG-1.0" ;
		:title = "California Underwater Glider Network - Line 90" ;
		:keywords = "AUVS > Autonomous Underwater Vehicles, Oceans > Ocean Pressure > Water Pressure, Oceans > Ocean Temperature > Water Temperature, Oceans > Salinity/Density > Conductivity, Oceans > Salinity/Density > Density, Oceans > Salinity/Density > Salinity" ;
		:keywords_vocabulary = "GCMD Science Keywords" ;
		:featureType = "trajectory" ;
		:id = "sp041-20191205T1757_R" ;
		:naming_authority = "edu.ucsd.spray" ;
		:history = "readsat - 2020-05-18T19:31:07Z, fixgps3 - 2020-05-18T19:31:07Z, calcvelsat - 2020-05-18T19:31:07Z, calox - 2021-02-26T11:39:46Z, addoxumolkg - 2021-02-26T11:39:46Z" ;
		:references = "Rudnick, D. L. (2016). Ocean research enabled by underwater gliders. Annual review of marine science, 8, 519-541, doi:10.1146/annurev-marine-122414-033913\n Rudnick, D. L., Davis, R. E., & Sherman, J. T. (2016). Spray Underwater Glider Operations. Journal of Atmospheric and Oceanic Technology, 33(6), 1113-1122, doi:10.1175/JTECH-D-15-0252.1\n Rudnick, D. L., Davis, R. E., Eriksen, C. C., Fratantoni, D. M., & Perry, M. J. (2004). Underwater gliders for ocean research. Marine Technology Society Journal, 38(2), 73-84, doi:10.4031/002533204787522703\n Sherman, J., Davis, R. E., Owens, W. B., & Valdes, J. (2001). The autonomous underwater glider \'Spray\'. IEEE Journal of oceanic Engineering, 26(4), 437-446, doi:10.1109/48.972076" ;
		:comment = "Dataset for demonstration purposes only. Original dataset truncated for the sake of simplicity" ;
		:processing_level = "Automatic quality control" ;
		:standard_name_vocabulary = "CF Standard Name Table v79" ;
		:date_created = "2022-08-17T06:54:43.077222" ;
		:creator_name = "Instrument Development Group" ;
		:creator_email = "idgdata@ucsd.edu" ;
		:creator_url = "http://spraydata.ucsd.edu" ;
		:creator_type = "group" ;
		:creator_institution = "University of California - San Diego; Scripps Institution of Oceanography" ;
		:institution = "Scripps Institution of Oceanography" ;
		:project = "California Underwater Glider Network" ;
		:publisher_name = "Instrument Development Group" ;
		:publisher_email = "idgdata@ucsd.edu" ;
		:publisher_url = "https://spraydata.ucsd.edu" ;
		:publisher_type = "group" ;
		:publisher_institution = "University of California - San Diego; Scripps Institution of Oceanography" ;
		:geospatial_bounds = "POLYGON ((-119.82769 32.50146, -119.821205 32.50548, -119.80175 32.51754, -119.82769 32.50146))" ;
		:geospatial_bounds_crs = "EPSG:4326" ;
		:geospatial_bounds_vertical_crs = "EPSG:5831" ;
		:geospatial_lat_min = 32.50146 ;
		:geospatial_lat_max = 32.51754 ;
		:geospatial_lon_min = -119.82769 ;
		:geospatial_lon_max = -119.80175 ;
		:geospatial_vertical_min = 1.54 ;
		:geospatial_vertical_max = 24.59 ;
		:geospatial_vertical_positive = "down" ;
		:geospatial_vertical_units = "m" ;
		:time_coverage_start = "2019-12-16T17:20:17Z" ;
		:time_coverage_end = "2019-12-16T17:23:13Z" ;
		:program = "GOMO, IOOS" ;
		:contributor_name = "Daniel Rudnick,Guilherme Castelao" ;
		:contributor_role = "Principal Investigator, Data Curator" ;
		:product_version = "v3" ;
		:platform = "Autonomous Underwater Vehicle" ;
		:instrument = "Seabird SBE 41CP" ;
		:metadata_link = "http://spraydata.ucsd.edu" ;
		:ctd_make_model = "Seabird SBE 41CP" ;
		:doi = "10.21238/S8SPRAY1618" ;
		:xglider_type = "trajectoryObs" ;
		:trajectory = "sp041-20191205T1757" ;
		:platform_vocabulary = "https://vocab.nerc.ac.uk/collection/L06/current/27/" ;
		:wmoid = "4801948" ;
		:internal_mission_identifier = "19C04101" ;
		:site = "CUGN line 90" ;
		:site_vocabulary = "TBD" ;
		:network = "California Underwater Glider Network" ;
		:contributor_email = "drudnick@ucsd.edu,castelao@ucsd.edu" ;
		:contributor_id = "0000-0002-2624-7074,0000-0002-6765-0708" ;
		:contributor_role_vocabulary = "https://orcid.org/" ;
		:agency = "Scripps Institution of Oceanography" ;
		:agency_role = "SDNPR004" ;
		:agency_role_vocabulary = "http://vocab.nerc.ac.uk/collection/C86/" ;
		:agency_id = "1390" ;
		:agency_id_vocabulary = "EDMO" ;
		:data_url = "https://spraydata.ucsd.edu/projects/CUGN/" ;
		:rtqc_method = "Spray - CoTeDe" ;
		:rtqc_method_doi = "10.21105/joss.02063" ;
		:web_link = "https://spraydata.ucsd.edu/projects/CUGN/" ;
		:mission = "19C04101" ;
		:date_modified = "2021-10-06T18:36:50.099674" ;
data:

 TRAJECTORY = "sp041-20191205T1757" ;

 PARAMETER = "PRES", "TEMP", "PSAL", "CHLA", "DOXY" ;

 TIME_GPS = 1576507260, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, 1576517403 ;

 TIME_GPS_QC = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _ ;

 LATITUDE_GPS = 32.51754, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, 32.50146 ;

 LATITUDE_GPS_QC = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _ ;

 LONGITUDE_GPS = -119.80175, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, -119.82769 ;

 LONGITUDE_GPS_QC = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _ ;

 PLATFORM = "sp041" ;

 PHASE = _, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, _ ;

 PHASE_QC = _, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, _ ;

 TIME = 1576507260, 1576516817, 1576516825, 1576516833, 1576516841, 
    1576516849, 1576516857, 1576516865, 1576516873, 1576516881, 1576516889, 
    1576516897, 1576516905, 1576516913, 1576516921, 1576516929, 1576516937, 
    1576516945, 1576516953, 1576516961, 1576516969, 1576516977, 1576516985, 
    1576516993, 1576517403 ;

 LATITUDE = 32.51754, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, 32.50146 ;

 LONGITUDE = -119.80175, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, -119.82769 ;

 PRES = _, 24.76, 23.68, 22.76, 21.72, 20.72, 19.68, 18.64, 17.48, 16.6, 
    15.52, 14.6, 13.44, 12.44, 11.4, 10.2, 8.44, 7.44, 6.28, 5.32, 4.36, 3.4, 
    2.32, 1.56, _ ;

 PRES_QC = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _ ;

 DEPTH = _, 24.5849769627501, 23.5126728256206, 22.5992241312562, 
    21.5666250478649, 20.5737364026879, 19.5411271039573, 18.5085125971717, 
    17.3567441183672, 16.4829843983173, 15.4106378268966, 14.4971529837432, 
    13.3453619368607, 12.3524334192887, 11.3197826520277, 10.1282560628289, 
    8.38067118597407, 7.38771858618288, 6.23588753584426, 5.28264314410755, 
    4.32939431287006, 3.37614104200687, 2.30372580539014, 1.5490598630261, _ ;

 TEMP = _, 15.505, 15.506, 15.505, 15.505, 15.506, 15.505, 15.505, 15.505, 
    15.504, 15.506, 15.504, 15.505, 15.508, 15.507, 15.509, 15.509, 15.51, 
    15.51, 15.511, 15.51, 15.511, 15.512, 15.512, _ ;

 TEMP_QC = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _ ;

 PSAL = _, 33.561, 33.561, 33.561, 33.561, 33.562, 33.561, 33.561, 33.561, 
    33.562, 33.561, 33.561, 33.561, 33.561, 33.561, 33.561, 33.561, 33.561, 
    33.56, 33.561, 33.56, 33.56, 33.559, 33.56, _ ;

 PSAL_QC = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _ ;

 DEPLOYMENT_TIME = 1575570735 ;

 DEPLOYMENT_LATITUDE = 32.9018 ;

 DEPLOYMENT_LONGITUDE = -117.299725 ;

 TELECOM_TYPE = "Iridium" ;

 TRACKING_SYSTEM = "GPS, ARGOS" ;

 N_MEASUREMENTS = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 
    17, 18, 19, 20, 21, 22, 23, 24 ;

 PLATFORM_TYPE = "Spray" ;

 PLATFORM_MODEL = "Spray" ;

 PLATFORM_MAKER = "Scripps Institution of Oceanography" ;

 PLATFORM_SERIAL_NUMBER = "0041" ;

 PLATFORM_CODE = "sp041" ;

 PLATFORM_DEPTH_RATING = 1000 ;

 WMO_IDENTIFIER = "4801948" ;

group: CTD {

  // group attributes:
  		:long_name = "Sea-Bird SBE 41CP CTD" ;
  		:type = "CTD" ;
  		:type_vocabulary = "https://vocab.nerc.ac.uk/collection/L05/current/130/" ;
  		:maker = "Sea-Bird Scientific" ;
  		:maker_vocabulary = "https://vocab.nerc.ac.uk/collection/L35/current/MAN0013/" ;
  		:model = "SBE 41CP CTD " ;
  		:model_vocabulary = "https://vocab.nerc.ac.uk/collection/L22/current/TOOL0669/" ;
  		:serial_number = "75" ;
  		:calibration_date = "2019-10-22T00:00:00Z" ;
  } // group CTD

group: OPTODE_DOXY {

  // group attributes:
  		:long_name = "Sea-Bird SBE 63 dissolved oxygen sensor" ;
  		:type = "OPTODE_DOXY" ;
  		:type_vocabulary = "https://vocab.nerc.ac.uk/collection/L05/current/351/" ;
  		:maker = "Seabird" ;
  		:maker_vocabulary = "https://vocab.nerc.ac.uk/collection/L35/current/MAN0013/" ;
  		:model = "Sea-Bird SBE 63 DO" ;
  		:model_identifier = "https://vocab.nerc.ac.uk/collection/L22/current/TOOL0739/" ;
  		:serial_number = "631776" ;
  		:calibration_date = "2019-11-22T00:00:00Z" ;
  } // group OPTODE_DOXY

group: FLUOROMETER_CHLA {
  dimensions:
  	N_MEASUREMENTS = 25 ;
  variables:
  	double CHLA(N_MEASUREMENTS) ;
  		CHLA:_FillValue = NaN ;
  		CHLA:long_name = "Chlorophyll-a concentration" ;
  		CHLA:standard_name = "mass_concentration_of_chlorophyll_a_in_sea_water" ;
  		CHLA:units = "mg m-3" ;
  		CHLA:ancillary_variables = "CHLA_QC" ;
  		CHLA:coverage_content_type = "physicalMeasurement" ;
  		CHLA:coordinates = "time lon lat depth" ;
  		CHLA:comment = "In-situ fluorometer with either manufacturer, laboratory or sample calibration applied" ;
  	byte CHLA_QC(N_MEASUREMENTS) ;
  		CHLA_QC:_FillValue = 0b ;
  		CHLA_QC:long_name = "quality flag" ;
  	int N_MEASUREMENTS(N_MEASUREMENTS) ;

  // group attributes:
  		:long_name = "Seapoint chlorophyll fluorometer" ;
  		:type = "FLUOROMETER_CHLA" ;
  		:type_vocabulary = "https://vocab.nerc.ac.uk/collection/L05/current/113/" ;
  		:maker = "SEAPOINT" ;
  		:maker_vocabulary = "https://vocab.nerc.ac.uk/collection/L35/current/MAN0177/" ;
  		:model = "Seapoint SCF" ;
  		:model_identifier = "http://vocab.nerc.ac.uk/collection/L22/current/TOOL0119/" ;
  		:serial_number = "S-5012" ;
  		:calibration_date = "2019-11-22T00:00:00Z" ;
  data:

   CHLA = _, 0.861, 0.909, 0.873, 0.867, 0.834, 0.864, 0.882, 0.855, 0.93, 
      0.819, 0.786, 0.807, 0.783, 0.741, 0.744, 0.609, 0.555, 0.573, 0.498, 
      0.471, 0.453, 0.444, 0.414, _ ;

   CHLA_QC = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
      _, _, _, _ ;

   N_MEASUREMENTS = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 
      17, 18, 19, 20, 21, 22, 23, 24 ;
  } // group FLUOROMETER_CHLA
}

netcdf sp041_20191205T1757 {
    dimensions:
        N_MEASUREMENTS = 25 ;
    variables:
        double LATITUDE_GPS(N_MEASUREMENTS) ;
            LATITUDE_GPS:long_name = "latitude of each GPS location" ;
            LATITUDE_GPS:standard_name = "latitude" ;
            LATITUDE_GPS:units = "degrees_north" ;
            LATITUDE_GPS:_FillValue = -9999.9 ;
            LATITUDE_GPS:valid_max = "90" ;
            LATITUDE_GPS:valid_min = "-90" ;
            LATITUDE_GPS:ancillary_variables = "LATITUDE_GPS_QC" ;
        double LONGITUDE_GPS(N_MEASUREMENTS) ;
            LONGITUDE_GPS:long_name = "longitude of each GPS location" ;
            LONGITUDE_GPS:standard_name = "longitude" ;
            LONGITUDE_GPS:units = "degrees_east" ;
            LONGITUDE_GPS:_FillValue = -9999.9 ;
            LONGITUDE_GPS:valid_max = "180" ;
            LONGITUDE_GPS:valid_min = "-180" ;
            LONGITUDE_GPS:ancillary_variables = "LONGITUDE_GPS_QC" ;
        double TIME_GPS(N_MEASUREMENTS) ;
            TIME_GPS:long_name = "time of each GPS location" ;
            TIME_GPS:calendar = "gregorian" ;
            TIME_GPS:units = "seconds since 1970-01-01T00:00:00Z" ;
            TIME_GPS:_FillValue = -1. ;
            TIME_GPS:valid_min = 1e9 ;
            TIME_GPS:valid_max = 4e9 ;
            TIME_GPS:ancillary_variables = "TIME_GPS_QC" ;
        double LATITUDE(N_MEASUREMENTS) ;
            LATITUDE:long_name = "latitude of each measurement and GPS location" ;
            LATITUDE:standard_name = "latitude" ;
            LATITUDE:units = "degrees_north" ;
            LATITUDE:_FillValue = -9999.9 ;
            LATITUDE:valid_min = "-90" ;
            LATITUDE:valid_max = "90" ;
            LATITUDE:ancillary_variables = "LATITUDE_GPS_QC"
            LATITUDE:interpolation_methodology = "TBD" ;
            LATITUDE:interpolation_methodology_vocabulary = "TBD" ;
            LATITUDE:interpolation_methodology_doi = "TBD" ;
        double LONGITUDE(N_MEASUREMENTS) ;
            LONGITUDE:long_name = "longitude of each measurements and GPS locations" ;
            LONGITUDE:standard_name = "longitude" ;
            LONGITUDE:units = "degrees_east" ;
            LONGITUDE:_FillValue = -9999.9 ;
            LONGITUDE:valid_min = "-180" ;
            LONGITUDE:valid_max = "180" ;
            LONGITUDE:ancillary_variables = "LONGITUDE_GPS_QC";
            LONGITUDE:interpolation_methodology = "TBD" ;
            LONGITUDE:interpolation_methodology_vocabulary = "TBD" ;
            LONGITUDE:interpolation_methodology_doi = "TBD" ;
        double TIME(N_MEASUREMENTS) ;
            TIME:long_name = "time of measurement and GPS location" ;
            TIME:calendar = "gregorian" ;
            TIME:units = "seconds since 1970-01-01T00:00:00Z" ;
            TIME:_FillValue = -1. ;
            TIME:valid_min = 1e9 ;
            TIME:valid_max = 4e9 ;
            TIME:interpolation_methodology = "TBD" ;
            TIME:interpolation_methodology_vocabulary = "TBD" ;
            TIME:interpolation_methodology_doi = "TBD" ;
        string TRAJECTORY ;
            TRAJECTORY:cf_role = "trajectory_id";
            TRAJECTORY:long_name = "trajectory name";
        string PLATFORM_MODEL ;
            PLATFORM_MODEL:long_name = "model of the glider" ;
            PLATFORM_MODEL:platform_model_vocabulary = "http://vocab.nerc.ac.uk/collection/B76/current/";
        string WMO_IDENTIFIER ;
            WMO_IDENTIFIER:long_name = "wmo id" ;
        double DEPLOYMENT_TIME ;
            DEPLOYMENT_TIME:long_name = "date of deployment" ;
            DEPLOYMENT_TIME:standard_name = "time" ;
            DEPLOYMENT_TIME:calendar = "gregorian" ;
            DEPLOYMENT_TIME:units = "seconds since 1970-01-01T00:00:00Z" ;
        double DEPLOYMENT_LATITUDE ;
            DEPLOYMENT_LATITUDE:long_name = "latitude of deployment" ;
            DEPLOYMENT_LATITUDE:standard_name = "latitude" ;
            DEPLOYMENT_LATITUDE:units = "degrees_north" ;
            DEPLOYMENT_LATITUDE:valid_max = "90" ;
            DEPLOYMENT_LATITUDE:valid_min = "-90" ;
        double DEPLOYMENT_LONGITUDE ;
            DEPLOYMENT_LONGITUDE:long_name = "longitude of deployment" ;
            DEPLOYMENT_LONGITUDE:standard_name = "longitude" ;
            DEPLOYMENT_LONGITUDE:units = "degrees_east" ;
            DEPLOYMENT_LONGITUDE:valid_max = "180" ;
            DEPLOYMENT_LONGITUDE:valid_min = "-180" ;
        float PRES(N_MEASUREMENTS) ;
            PRES:long_name = "Pressure" ;
            PRES:standard_name = "sea_water_pressure" ;
            PRES:vocabulary = "http://vocab.nerc.ac.uk/collection/OG1/current/PRES/";
            PRES:_FillValue = -9999.9 ;
            PRES:units = "dbar" ;
            PRES:ancillary_variables = "PRES_QC" ;
            PRES:coordinates = "LATITUDE, LONGITUDE, DEPTH, TIME" ;
        float DEPTH(N_MEASUREMENTS) ;
            DEPTH:long_name = "Depth" ;
            DEPTH:standard_name = "depth" ;
            DEPTH:vocabulary = "http://vocab.nerc.ac.uk/collection/OG1/current/DEPTH/";
            DEPTH:_FillValue = NaN ;
            DEPTH:units = "m" ;
            DEPTH:ancillary_variables = "DEPTH_QC" ;
            DEPTH:coordinates = "LATITUDE, LONGITUDE, DEPTH, TIME" ;
        float TEMP(N_MEASUREMENTS) ;
            TEMP:long_name = "Sea Water Temperature" ;
            TEMP:standard_name = "sea_water_temperature" ;
            TEMP:vocabulary = "http://vocab.nerc.ac.uk/collection/OG1/current/TEMP/";
            TEMP:_FillValue = -9999.9 ;
            TEMP:units = "Celsius" ;
            TEMP:ancillary_variables = "TEMP_QC" ;
            TEMP:coordinates = "LATITUDE, LONGITUDE, DEPTH, TIME" ;
        float PSAL(N_MEASUREMENTS) ;
            PSAL:long_name = "Sea Water Salinity" ;
            PSAL:standard_name = "sea_water_practical_salinity" ;
            PSAL:vocabulary = "http://vocab.nerc.ac.uk/collection/OG1/current/PSAL/";
            PSAL:_FillValue = NaN ;
            PSAL:units = "1" ;
            PSAL:ancillary_variables = "PSAL_QC" ;
            PSAL:coordinates = "LATITUDE, LONGITUDE, DEPTH, TIME" ;
        float CHLA(N_MEASUREMENTS) ;
            CHLA:long_name = "Chlorophyll-a concentration" ;
            CHLA:standard_name = "mass_concentration_of_chlorophyll_a_in_sea_water" ;
            CHLA:vocabulary = "http://vocab.nerc.ac.uk/collection/OG1/current/CHLA/";
            CHLA:_FillValue = NaN ;
            CHLA:units = "mg m-3" ;
            CHLA:ancillary_variables = "CHLA_QC" ;
            CHLA:coordinates = "LATITUDE, LONGITUDE, DEPTH, TIME" ;
        float DOXY(N_MEASUREMENTS) ;
            DOXY:long_name = "Dissolved oxygen" ;
            DOXY:standard_name = "moles_of_oxygen_per_unit_mass_in_sea_water" ;
            DOXY:vocabulary = "http://vocab.nerc.ac.uk/collection/OG1/current/DOXY/";
            DOXY:_FillValue = NaN ;
            DOXY:units = "micromol kg-1" ;
            DOXY:ancillary_variables = "DOXY_QC" ;
            DOXY:coordinates = "LATITUDE, LONGITUDE, DEPTH, TIME" ;
    
    // global attributes:
            :title = "California Underwater Glider Network - Line 90" ;
            :platform = "sub-surface gliders" ;
            :platform_vocabulary = "https://vocab.nerc.ac.uk/collection/L06/current/27/" ;
            :id = "sp041_20191205T1757_R" ;
            :contributor_name = "Daniel Rudnick" ;
            :contributor_email = "drudnick@ucsd.edu" ;
            :contributor_role = "Principal Investigator" ;
            :contributor_role_vocabulary = "http://vocab.nerc.ac.uk/collection/W08/current/CONT0004/" ;
            :agency = "Scripps Institution of Oceanography" ;
            :agency_role = "programme operation responsibility" ;
            :agency_role_vocabulary = "http://vocab.nerc.ac.uk/collection/C86/current/SDNPR002/" ;
            :data_url = "https://spraydata.ucsd.edu/projects/CUGN/" ;
            :rtqc_method = "Spray - CoTeDe" ;
            :rtqc_method_doi = "10.21105/joss.02063" ;
            :date_created = "2021-04-10T01:14:44" ;
            :featureType = "trajectory" ;
            :Conventions = "CF-1.8, ACDD-1.3, OG-1.0" ;

    data:
    
     TRAJECTORY = "sp041_20191205T1757" ;
    
     PARAMETER = "PRES", "TEMP", "PSAL", "CHLA", "DOXY" ;
    
     TIME_GPS = 1576507260, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
        _, _, _, _, _, 1576517403 ;
    
     LATITUDE_GPS = 32.51754, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
        _, _, _, _, _, _, 32.50146 ;
    
     LONGITUDE_GPS = -119.80175, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
        _, _, _, _, _, _, _, -119.82769 ;
    
     TIME = 1576507260, 1576516817, 1576516825, 1576516833, 1576516841, 
        1576516849, 1576516857, 1576516865, 1576516873, 1576516881, 1576516889, 
        1576516897, 1576516905, 1576516913, 1576516921, 1576516929, 1576516937, 
        1576516945, 1576516953, 1576516961, 1576516969, 1576516977, 1576516985, 
        1576516993, 1576517403 ;
    
     LATITUDE = 32.51754, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
        _, _, _, _, _, 32.50146 ;
    
     LONGITUDE = -119.80175, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
        _, _, _, _, _, _, -119.82769 ;
    
     PRES = _, 24.76, 23.68, 22.76, 21.72, 20.72, 19.68, 18.64, 17.48, 16.6, 
        15.52, 14.6, 13.44, 12.44, 11.4, 10.2, 8.44, 7.44, 6.28, 5.32, 4.36, 3.4, 
        2.32, 1.56, _ ;
    
     DEPTH = _, 24.5849769627501, 23.5126728256206, 22.5992241312562, 
        21.5666250478649, 20.5737364026879, 19.5411271039573, 18.5085125971717, 
        17.3567441183672, 16.4829843983173, 15.4106378268966, 14.4971529837432, 
        13.3453619368607, 12.3524334192887, 11.3197826520277, 10.1282560628289, 
        8.38067118597407, 7.38771858618288, 6.23588753584426, 5.28264314410755, 
        4.32939431287006, 3.37614104200687, 2.30372580539014, 1.5490598630261, _ ;
    
     TEMP = _, 15.505, 15.506, 15.505, 15.505, 15.506, 15.505, 15.505, 15.505, 
        15.504, 15.506, 15.504, 15.505, 15.508, 15.507, 15.509, 15.509, 15.51, 
        15.51, 15.511, 15.51, 15.511, 15.512, 15.512, _ ;
    
     PSAL = _, 33.561, 33.561, 33.561, 33.561, 33.562, 33.561, 33.561, 33.561, 
        33.562, 33.561, 33.561, 33.561, 33.561, 33.561, 33.561, 33.561, 33.561, 
        33.56, 33.561, 33.56, 33.56, 33.559, 33.56, _ ;
    
     CHLA = _, 0.861, 0.909, 0.873, 0.867, 0.834, 0.864, 0.882, 0.855, 0.93, 
        0.819, 0.786, 0.807, 0.783, 0.741, 0.744, 0.609, 0.555, 0.573, 0.498, 
        0.471, 0.453, 0.444, 0.414, _ ;
    
     DOXY = _, 240.699500381006, 240.728111146589, 240.75690836507, 
        240.710612669174, 240.922144300944, 240.655413148225, 240.720151525978, 
        240.635340339479, 240.700230807224, 240.76636985969, 240.831706998232, 
        240.7111499353, 240.664998530651, 240.915858055632, 240.904784287258, 
        241.074164770971, 240.990908679491, 241.093556991221, 241.119569863555, 
        241.297597492548, 241.067163480339, 241.244566377113, 241.199209516033, _ ;
    
     DEPLOYMENT_TIME = 1575570735.0 ;
    
     DEPLOYMENT_LATITUDE = 32.9018 ;
    
     DEPLOYMENT_LONGITUDE = -117.29972500000001 ;
    
     PLATFORM_MODEL = "Spray" ;
    
     WMO_IDENTIFIER = "4801948" ;
    }

netcdf file:/Users/sevadjian/projects/og-netcdf/2022_11_test/og-10-CF18-for-cdl.nc {
  dimensions:
    N_PARAMS = 3;
    PARAM_STRLEN = 16;
    N_MEASUREMENTS = 4564;
    TRAJ_STRLEN = 19;
  variables:
    char TRAJECTORY(TRAJ_STRLEN=19);
      :cf_role = "trajectory_id";

    double TIME(N_MEASUREMENTS=4564);
      :axis = "T";
      :units = "seconds since 1970-01-01 00:00:00 UTC";
      :calendar = "julian";
      :standard_name = "time";
      :long_name = "Time";

    double LATITUDE(N_MEASUREMENTS=4564);
      :long_name = "Latitude";
      :standard_name = "latitude";
      :axis = "Y";
      :units = "degrees_north";

    double LONGITUDE(N_MEASUREMENTS=4564);
      :standard_name = "longitude";
      :axis = "X";
      :units = "degrees_east";
      :long_name = "Longitude";

    float DEPTH(N_MEASUREMENTS=4564);
      :positive = "down";
      :long_name = "Depth";
      :standard_name = "depth";
      :units = "m";
      :axis = "Z";

    double CHLA(N_MEASUREMENTS=4564);
      :_FillValue = -9999.0; // double
      :coordinates = "TIME LATITUDE LONGITUDE DEPTH";
      :standard_name = "mass_concentration_of_chlorophyll_a_in_sea_water";
      :long_name = "Chlorophyll-a concentration";
      :units = "mg m-3";
      :vocabulary = "https://vocab.nerc.ac.uk/collection/OG1/current/";
      :ancillary_variables = "CHLA_INSTRUMENT";

    float DENSITY(N_MEASUREMENTS=4564);
      :vocabulary = "https://vocab.nerc.ac.uk/collection/OG1/current/";
      :standard_name = "sea_water_density";
      :long_name = "Sea Water Density";
      :units = "kg m-3";
      :_FillValue = -9999.0f; // float
      :coordinates = "TIME LATITUDE LONGITUDE DEPTH";

    double DOXY(N_MEASUREMENTS=4564);
      :_FillValue = -9999.0; // double
      :coordinates = "TIME LATITUDE LONGITUDE DEPTH";
      :standard_name = "moles_of_oxygen_per_unit_mass_in_sea_water";
      :long_name = "Dissolved oxygen";
      :units = "micromol kg-1";
      :vocabulary = "https://vocab.nerc.ac.uk/collection/OG1/current/";
      :ancillary_variables = "DOXY_QC DOXY_INSTRUMENT";

    char PARAMETERS(N_PARAMS=3, PARAM_STRLEN=16);

    byte DOXY_QC(N_MEASUREMENTS=4564);
      :coordinates = "TIME LATITUDE LONGITUDE DEPTH";
      :long_name = "dissolved_oxygen Quality Flag";

    int CHLA_INSTRUMENT(N_MEASUREMENTS=4564);
      :long_name = "dissolved_oxygen Quality Flag";
      :vocabulary = "https://docs.google.com/document/d/1dN90xkw9oCbLs0sPPhOmszdOjLpwcqxiK5mjeZP7abA/edit";
      :make_model = "ECO_FL";

    int DOXY_INSTRUMENT(N_MEASUREMENTS=4564);
      :vocabulary = "https://docs.google.com/document/d/1dN90xkw9oCbLs0sPPhOmszdOjLpwcqxiK5mjeZP7abA/edit";
      :make_model = "SEABIRD_SBE43F_IDO";
      :long_name = "Dissolved Oxygen Instrument";

  // global attributes:
  :acknowledgement = "Funded by National Oceanic and Atmospheric Administration (NOAA): Global Ocean Monitoring and Observing (GOMO) Program and Integrated Ocean Observing System. Supported by Instrument Development Group - Scripps Institution of Oceanography";
  :contributor_name = "Daniel Rudnick, Jennifer Sevadjian";
  :contributor_role = "principalInvestigator, resourceProvider";
  :contributor_role_vocabulary = "https://vocab.nerc.ac.uk/collection/G04/current";
  :Conventions = "Unidata Dataset Discovery v1.0, COARDS, CF-1.8";
  :creator_email = "idgdata@ucsd.edu";
  :creator_institution = "Scripps Institution of Oceanography";
  :creator_name = "Instrument Development Group";
  :creator_type = "group";
  :creator_url = "https://spraydata.ucsd.edu";
  :date_created = "2023-01-24T16:20:56.349455";
  :date_issued = "2023-01-24T16:21:36.025291";
  :date_modified = "2023-01-24T16:21:24.465881";
  :doi = "10.21238/S8SPRAY1618";
  :Easternmost_Easting = -124.49495; // double
  :featureType = "trajectory";
  :format_version = "IOOS_Glider_NetCDF_v3.0.nc";
  :geospatial_bounds = "POLYGON ((-123.2773 38.3228, -123.278675 38.32355, -123.2828 38.3258, -123.2773 38.3228))";
  :geospatial_bounds_crs = "EPSG:4326";
  :geospatial_bounds_vertical_crs = "EPSG:5831";
  :geospatial_lat_max = 37.96675; // double
  :geospatial_lat_min = 37.43285; // double
  :geospatial_lat_units = "degrees_north";
  :geospatial_lon_max = -124.49495; // double
  :geospatial_lon_min = -125.99015; // double
  :geospatial_lon_units = "degrees_east";
  :geospatial_vertical_max = 502.2962f; // float
  :geospatial_vertical_min = 0.5955232f; // float
  :geospatial_vertical_positive = "down";
  :geospatial_vertical_units = "m";
  :gts_ingest = "true";
  :history = "readsat - 2023-01-24T08:20:39Z, fixgps3 - 2023-01-24T08:20:39Z, calcvelsat - 2023-01-24T08:20:39Z, autoqcctd - 2023-01-24T08:20:39Z, calox - 2023-01-24T08:20:40Z, calfchl - 2023-01-24T08:20:42Z, adpsat - 2023-01-24T08:20:52Z\n2023-04-24T16:53:57Z (local files)\n2023-04-24T16:53:57Z https://gliders.ioos.us/erddap/tabledap/sp011-20221014T1612.ncCF?&time%3E=1667088000.0&time%3C=1667692800.0";
  :id = "sp011-20221014T1612";
  :infoUrl = "https://gliders.ioos.us/erddap/";
  :institution = "Scripps Institution of Oceanography";
  :ioos_dac_checksum = "d4db73cb25d1345fca338bd5fc6f8db3";
  :ioos_dac_completed = "True";
  :keywords = "AUVS > Autonomous Underwater Vehicles, Earth Science > Oceans > Ocean Pressure > Water Pressure, Earth Science > Oceans > Ocean Temperature > Water Temperature, Earth Science > Oceans > Salinity/Density > Conductivity, Earth Science > Oceans > Salinity/Density > Density, Earth Science > Oceans > Salinity/Density > Salinity, glider, In Situ Ocean-based platforms > Seaglider, Slocum, Spray, trajectory, underwater glider, water, wmo";
  :keywords_vocabulary = "GCMD Science Keywords";
  :license = "Creative Commons Attribution 4.0 International Public License (https://creativecommons.org/licenses/by/4.0/)";
  :Metadata_Conventions = "Unidata Dataset Discovery v1.0, COARDS, CF-1.6";
  :metadata_link = "https://spraydata.ucsd.edu";
  :naming_authority = "edu.ucsd.idg";
  :network = "OceanGliders > BOON > Northeast Pacific Ocean > California Underwater Glider Network, California Underwater Glider Network (CUGN), IOOS";
  :Northernmost_Northing = 37.96675; // double
  :platform = "sp011";
  :platform_institution = "Scripps Institution of Oceanography";
  :platform_type = "Spray Glider";
  :processing_level = "Level 2 - Real-time automatic quality control has been applied. Data quality flags have been added. See the infoUrl for more information about data processing for this data stream as well as information about available data products with additional processing applied.";
  :product_version = "v3";
  :project = "California Underwater Glider Network (CUGN)";
  :publisher_email = "idgdata@ucsd.edu";
  :publisher_institution = "University of California - San Diego; Scripps Institution of Oceanography";
  :publisher_name = "Instrument Development Group";
  :publisher_type = "group";
  :publisher_url = "https://spraydata.ucsd.edu";
  :references = "Rudnick, D. L. (2016). Ocean research enabled by underwater gliders. Annual review of marine science, 8, 519-541, doi:10.1146/annurev-marine-122414-033913\n Rudnick, D. L., Davis, R. E., & Sherman, J. T. (2016). Spray Underwater Glider Operations. Journal of Atmospheric and Oceanic Technology, 33(6), 1113-1122, doi:10.1175/JTECH-D-15-0252.1\n Rudnick, D. L., Davis, R. E., Eriksen, C. C., Fratantoni, D. M., & Perry, M. J. (2004). Underwater gliders for ocean research. Marine Technology Society Journal, 38(2), 73-84, doi:10.4031/002533204787522703\n Sherman, J., Davis, R. E., Owens, W. B., & Valdes, J. (2001). The autonomous underwater glider \'Spray\'. IEEE Journal of oceanic Engineering, 26(4), 437-446, doi:10.1109/48.972076";
  :sea_name = "Coastal Waters of California";
  :site = "CUGN Line 56";
  :source = "Observational data from a profiling underwater glider.";
  :sourceUrl = "(local files)";
  :Southernmost_Northing = 37.43285; // double
  :standard_name_vocabulary = "CF Standard Name Table v75";
  :subsetVariables = "wmo_id,trajectory,profile_id,time,latitude,longitude";
  :summary = "The overarching goal of the California Underwater Glider Network is to sustain baseline observations of climate variability off the coast of California. The technical approach is to deploy autonomous underwater gliders in a network to provide real-time data.\nThe CUGN uses Spray underwater gliders making repeated dives from the surface to 500 m and back, repeating the cycle every 3 hours, and traveling 3 km in the horizontal during that time. The CUGN includes gliders on three of the traditional cross-shore CalCOFI lines: line 66.7 off Monterey Bay, line 80 off Point Conception, and line 90 off Dana Point.\n The glider missions typically last about 100 days, and cover over 2000 km, thus providing 4-6 sections on lines extending 300-500 km offshore. Since 2005 the CUGN has covered 200,000 km over ground in 28 glider-years, while doing 90,000 dives.";
  :time_coverage_end = "2022-11-05T22:31:30Z";
  :time_coverage_start = "2022-10-30T00:19:30Z";
  :title = "sp011-20221014T1612";
  :trajectory = "sp011-20221014T1612";
  :Westernmost_Easting = -125.99015; // double
  :xglider_type = "profileObs";
  :cdm_data_type = "Trajectory";

  data:
    TRAJECTORY =   "sp011-20221014T1612"
    TIME = 
      {1.667082061E9, 1.667087871E9, 1.667087918E9, 1.667087966E9, 1.667088014E9, 1.667088062E9, 1.66708811E9, 1.667088158E9, 1.667088206E9, 1.667088254E9, 1.667088302E9, 1.66708835E9, 1.667088398E9, 1.667088446E9, 1.667088494E9, 1.667088542E9, 1.66708859E9, 1.667088638E9, 1.667088686E9, 1.667088734E9, 1.667088782E9, 1.66708883E9, 1.667088878E9, 1.667088926E9, 1.667088974E9, 1.667089022E9, 1.66708907E9, 1.667089118E9, 1.667089166E9, 1.667089214E9, 1.667089262E9, 1.66708931E9, 1.667089358E9, 1.667089406E9, 1.667089454E9, 1.667089502E9, 1.66708955E9, 1.667089598E9, 1.667089646E9, 1.667089694E9, 1.667089742E9, 1.66708979E9, 1.667089838E9, 1.667089886E9, 1.667089934E9, 1.667089982E9, 1.66709003E9, 1.667090078E9, 1.667090126E9, 1.667090174E9, 1.667090222E9, 1.66709027E9, 1.667090318E9, 1.667090366E9, 1.667090414E9, 1.667090462E9, 1.66709051E9, 1.667090558E9, 1.667090606E9, 1.667090654E9, 1.667090702E9, 1.66709075E9, 1.667090798E9, 1.667090846E9, 1.667090894E9, 1.667090942E9, 1.66709099E9, 1.667091038E9, 1.667091086E9, 1.667091134E9, 1.667091182E9, 1.66709123E9, 1.66709154E9, 1.66709172E9, 1.667097482E9, 1.66709753E9, 1.667097578E9, 1.667097626E9, 1.667097674E9, 1.667097722E9, 1.66709777E9, 1.667097818E9, 1.667097866E9, 1.667097914E9, 1.667097962E9, 1.66709801E9, 1.667098058E9, 1.667098106E9, 1.667098154E9, 1.667098202E9, 1.66709825E9, 1.667098298E9, 1.667098346E9, 1.667098394E9, 1.667098442E9, 1.66709849E9, 1.667098538E9, 1.667098586E9, 1.667098634E9, 1.667098682E9, 1.66709873E9, 1.667098778E9, 1.667098826E9, 1.667098874E9, 1.667098922E9, 1.66709897E9, 1.667099018E9, 1.667099066E9, 1.667099114E9, 1.667099162E9, 1.66709921E9, 1.667099258E9, 1.667099306E9, 1.667099354E9, 1.667099402E9, 1.66709945E9, 1.667099498E9, 1.667099546E9, 1.667099594E9, 1.667099642E9, 1.66709969E9, 1.667099738E9, 1.667099786E9, 1.667099834E9, 1.667099882E9, 1.66709993E9, 1.667099978E9, 1.667100026E9, 1.667100074E9, 1.667100122E9, 1.66710017E9, 1.667100218E9, 1.667100266E9, 1.667100314E9, 1.667100362E9, 1.66710041E9, 1.667100458E9, 1.667100506E9, 1.667100554E9, 1.667100602E9, 1.66710065E9, 1.66710096E9, 1.66710114E9, 1.667106857E9, 1.667106905E9, 1.667106953E9, 1.667107001E9, 1.667107049E9, 1.667107097E9, 1.667107145E9, 1.667107193E9, 1.667107241E9, 1.667107289E9, 1.667107337E9, 1.667107385E9, 1.667107433E9, 1.667107481E9, 1.667107529E9, 1.667107577E9, 1.667107625E9, 1.667107673E9, 1.667107721E9, 1.667107769E9, 1.667107817E9, 1.667107865E9, 1.667107913E9, 1.667107961E9, 1.667108009E9, 1.667108057E9, 1.667108105E9, 1.667108153E9, 1.667108201E9, 1.667108249E9, 1.667108297E9, 1.667108345E9, 1.667108393E9, 1.667108441E9, 1.667108489E9, 1.667108537E9, 1.667108585E9, 1.667108633E9, 1.667108681E9, 1.667108729E9, 1.667108777E9, 1.667108825E9, 1.667108873E9, 1.667108921E9, 1.667108969E9, 1.667109017E9, 1.667109065E9, 1.667109113E9, 1.667109161E9, 1.667109209E9, 1.667109257E9, 1.667109305E9, 1.667109353E9, 1.667109401E9, 1.667109449E9, 1.667109497E9, 1.667109545E9, 1.667109593E9, 1.667109641E9, 1.667109689E9, 1.667109737E9, 1.667109785E9, 1.667109833E9, 1.667109881E9, 1.667109929E9, 1.667109977E9, 1.667110025E9, 1.667110073E9, 1.667110121E9, 1.667110169E9, 1.6671105E9, 1.66711068E9, 1.667116457E9, 1.667116505E9, 1.667116553E9, 1.667116601E9, 1.667116649E9, 1.667116697E9, 1.667116745E9, 1.667116793E9, 1.667116841E9, 1.667116889E9, 1.667116937E9, 1.667116985E9, 1.667117033E9, 1.667117081E9, 1.667117129E9, 1.667117177E9, 1.667117225E9, 1.667117273E9, 1.667117321E9, 1.667117369E9, 1.667117417E9, 1.667117465E9, 1.667117513E9, 1.667117561E9, 1.667117609E9, 1.667117657E9, 1.667117705E9, 1.667117753E9, 1.667117801E9, 1.667117849E9, 1.667117897E9, 1.667117945E9, 1.667117993E9, 1.667118041E9, 1.667118089E9, 1.667118137E9, 1.667118185E9, 1.667118233E9, 1.667118281E9, 1.667118329E9, 1.667118377E9, 1.667118425E9, 1.667118473E9, 1.667118521E9, 1.667118569E9, 1.667118617E9, 1.667118665E9, 1.667118713E9, 1.667118761E9, 1.667118809E9, 1.667118857E9, 1.667118905E9, 1.667118953E9, 1.667119001E9, 1.667119049E9, 1.667119097E9, 1.667119145E9, 1.667119193E9, 1.667119241E9, 1.667119289E9, 1.667119337E9, 1.667119385E9, 1.667119433E9, 1.667119481E9, 1.667119529E9, 1.6671198E9, 1.66711998E9, 1.667125544E9, 1.667125592E9, 1.66712564E9, 1.667125688E9, 1.667125736E9, 1.667125784E9, 1.667125832E9, 1.66712588E9, 1.667125928E9, 1.667125976E9, 1.667126024E9, 1.667126072E9, 1.66712612E9, 1.667126168E9, 1.667126216E9, 1.667126264E9, 1.667126312E9, 1.66712636E9, 1.667126408E9, 1.667126456E9, 1.667126504E9, 1.667126552E9, 1.6671266E9, 1.667126648E9, 1.667126696E9, 1.667126744E9, 1.667126792E9, 1.66712684E9, 1.667126888E9, 1.667126936E9, 1.667126984E9, 1.667127032E9, 1.66712708E9, 1.667127128E9, 1.667127176E9, 1.667127224E9, 1.667127272E9, 1.66712732E9, 1.667127368E9, 1.667127416E9, 1.667127464E9, 1.667127512E9, 1.66712756E9, 1.667127608E9, 1.667127656E9, 1.667127704E9, 1.667127752E9, 1.6671278E9, 1.667127848E9, 1.667127896E9, 1.667127944E9, 1.667127992E9, 1.66712804E9, 1.667128088E9, 1.667128136E9, 1.667128184E9, 1.667128232E9, 1.66712828E9, 1.667128328E9, 1.667128376E9, 1.667128424E9, 1.667128472E9, 1.66712852E9, 1.667128568E9, 1.667128616E9, 1.667128664E9, 1.667128712E9, 1.66712876E9, 1.6671291E9, 1.66712928E9, 1.667134992E9, 1.66713504E9, 1.667135088E9, 1.667135136E9, 1.667135184E9, 1.667135232E9, 1.66713528E9, 1.667135328E9, 1.667135376E9, 1.667135424E9, 1.667135472E9, 1.66713552E9, 1.667135568E9, 1.667135616E9, 1.667135664E9, 1.667135712E9, 1.66713576E9, 1.667135808E9, 1.667135856E9, 1.667135904E9, 1.667135952E9, 1.667136E9, 1.667136048E9, 1.667136096E9, 1.667136144E9, 1.667136192E9, 1.66713624E9, 1.667136288E9, 1.667136336E9, 1.667136384E9, 1.667136432E9, 1.66713648E9, 1.667136528E9, 1.667136576E9, 1.667136624E9, 1.667136672E9, 1.66713672E9, 1.667136768E9, 1.667136816E9, 1.667136864E9, 1.667136912E9, 1.66713696E9, 1.667137008E9, 1.667137056E9, 1.667137104E9, 1.667137152E9, 1.6671372E9, 1.667137248E9, 1.667137296E9, 1.667137344E9, 1.667137392E9, 1.66713744E9, 1.667137488E9, 1.667137536E9, 1.667137584E9, 1.667137632E9, 1.66713768E9, 1.667137728E9, 1.667137776E9, 1.667137824E9, 1.667137872E9, 1.66713792E9, 1.667137968E9, 1.667138016E9, 1.667138064E9, 1.667138112E9, 1.66713816E9, 1.667138208E9, 1.667138256E9, 1.667138304E9, 1.667138352E9, 1.6671384E9, 1.66713876E9, 1.66713906E9, 1.667144845E9, 1.667144893E9, 1.667144941E9, 1.667144989E9, 1.667145037E9, 1.667145085E9, 1.667145133E9, 1.667145181E9, 1.667145229E9, 1.667145277E9, 1.667145325E9, 1.667145373E9, 1.667145421E9, 1.667145469E9, 1.667145517E9, 1.667145565E9, 1.667145613E9, 1.667145661E9, 1.667145709E9, 1.667145757E9, 1.667145805E9, 1.667145853E9, 1.667145901E9, 1.667145949E9, 1.667145997E9, 1.667146045E9, 1.667146093E9, 1.667146141E9, 1.667146189E9, 1.667146237E9, 1.667146285E9, 1.667146333E9, 1.667146381E9, 1.667146429E9, 1.667146477E9, 1.667146525E9, 1.667146573E9, 1.667146621E9, 1.667146669E9, 1.667146717E9, 1.667146765E9, 1.667146813E9, 1.667146861E9, 1.667146909E9, 1.667146957E9, 1.667147005E9, 1.667147053E9, 1.667147101E9, 1.667147149E9, 1.667147197E9, 1.667147245E9, 1.667147293E9, 1.667147341E9, 1.667147389E9, 1.667147437E9, 1.667147485E9, 1.667147533E9, 1.667147581E9, 1.667147629E9, 1.667147677E9, 1.667147725E9, 1.667147773E9, 1.667147821E9, 1.667147869E9, 1.667147917E9, 1.667147965E9, 1.667148013E9, 1.667148061E9, 1.667148109E9, 1.66714842E9, 1.6671486E9, 1.667154155E9, 1.667154203E9, 1.667154251E9, 1.667154299E9, 1.667154347E9, 1.667154395E9, 1.667154443E9, 1.667154491E9, 1.667154539E9, 1.667154587E9, 1.667154635E9, 1.667154683E9, 1.667154731E9, 1.667154779E9, 1.667154827E9, 1.667154875E9, 1.667154923E9, 1.667154971E9, 1.667155019E9, 1.667155067E9, 1.667155115E9, 1.667155163E9, 1.667155211E9, 1.667155259E9, 1.667155307E9, 1.667155355E9, 1.667155403E9, 1.667155451E9, 1.667155499E9, 1.667155547E9, 1.667155595E9, 1.667155643E9, 1.667155691E9, 1.667155739E9, 1.667155787E9, 1.667155835E9, 1.667155883E9, 1.667155931E9, 1.667155979E9, 1.667156027E9, 1.667156075E9, 1.667156123E9, 1.667156171E9, 1.667156219E9, 1.667156267E9, 1.667156315E9, 1.667156363E9, 1.667156411E9, 1.667156459E9, 1.667156507E9, 1.667156555E9, 1.667156603E9, 1.667156651E9, 1.667156699E9, 1.667156747E9, 1.667156795E9, 1.667156843E9, 1.667156891E9, 1.667156939E9, 1.667156987E9, 1.667157035E9, 1.667157083E9, 1.667157131E9, 1.667157179E9, 1.667157227E9, 1.667157275E9, 1.667157323E9, 1.667157371E9, 1.667157419E9, 1.66715772E9, 1.6671579E9, 1.667163741E9, 1.667163789E9, 1.667163837E9, 1.667163885E9, 1.667163933E9, 1.667163981E9, 1.667164029E9, 1.667164077E9, 1.667164125E9, 1.667164173E9, 1.667164221E9, 1.667164269E9, 1.667164317E9, 1.667164365E9, 1.667164413E9, 1.667164461E9, 1.667164509E9, 1.667164557E9, 1.667164605E9, 1.667164653E9, 1.667164701E9, 1.667164749E9, 1.667164797E9, 1.667164845E9, 1.667164893E9, 1.667164941E9, 1.667164989E9, 1.667165037E9, 1.667165085E9, 1.667165133E9, 1.667165181E9, 1.667165229E9, 1.667165277E9, 1.667165325E9, 1.667165373E9, 1.667165421E9, 1.667165469E9, 1.667165517E9, 1.667165565E9, 1.667165613E9, 1.667165661E9, 1.667165709E9, 1.667165757E9, 1.667165805E9, 1.667165853E9, 1.667165901E9, 1.667165949E9, 1.667165997E9, 1.667166045E9, 1.667166093E9, 1.667166141E9, 1.667166189E9, 1.667166237E9, 1.667166285E9, 1.667166333E9, 1.667166381E9, 1.667166429E9, 1.667166477E9, 1.667166525E9, 1.667166573E9, 1.667166621E9, 1.667166669E9, 1.667166717E9, 1.667166765E9, 1.667166813E9, 1.667166861E9, 1.667166909E9, 1.667166957E9, 1.667167005E9, 1.667167053E9, 1.667167101E9, 1.667167149E9, 1.6671675E9, 1.66716768E9, 1.66717351E9, 1.667173558E9, 1.667173606E9, 1.667173654E9, 1.667173702E9, 1.66717375E9, 1.667173798E9, 1.667173846E9, 1.667173894E9, 1.667173942E9, 1.66717399E9, 1.667174038E9, 1.667174086E9, 1.667174134E9, 1.667174182E9, 1.66717423E9, 1.667174278E9, 1.667174326E9, 1.667174374E9, 1.667174422E9, 1.66717447E9, 1.667174518E9, 1.667174566E9, 1.667174614E9, 1.667174662E9, 1.66717471E9, 1.667174758E9, 1.667174806E9, 1.667174854E9, 1.667174902E9, 1.66717495E9, 1.667174998E9, 1.667175046E9, 1.667175094E9, 1.667175142E9, 1.66717519E9, 1.667175238E9, 1.667175286E9, 1.667175334E9, 1.667175382E9, 1.66717543E9, 1.667175478E9, 1.667175526E9, 1.667175574E9, 1.667175622E9, 1.66717567E9, 1.667175718E9, 1.667175766E9, 1.667175814E9, 1.667175862E9, 1.66717591E9, 1.667175958E9, 1.667176006E9, 1.667176054E9, 1.667176102E9, 1.66717615E9, 1.667176198E9, 1.667176246E9, 1.667176294E9, 1.667176342E9, 1.66717639E9, 1.667176438E9, 1.667176486E9, 1.667176534E9, 1.667176582E9, 1.66717663E9, 1.66717692E9, 1.6671771E9, 1.667182933E9, 1.667182981E9, 1.667183029E9, 1.667183077E9, 1.667183125E9, 1.667183173E9, 1.667183221E9, 1.667183269E9, 1.667183317E9, 1.667183365E9, 1.667183413E9, 1.667183461E9, 1.667183509E9, 1.667183557E9, 1.667183605E9, 1.667183653E9, 1.667183701E9, 1.667183749E9, 1.667183797E9, 1.667183845E9, 1.667183893E9, 1.667183941E9, 1.667183989E9, 1.667184037E9, 1.667184085E9, 1.667184133E9, 1.667184181E9, 1.667184229E9, 1.667184277E9, 1.667184325E9, 1.667184373E9, 1.667184421E9, 1.667184469E9, 1.667184517E9, 1.667184565E9, 1.667184613E9, 1.667184661E9, 1.667184709E9, 1.667184757E9, 1.667184805E9, 1.667184853E9, 1.667184901E9, 1.667184949E9, 1.667184997E9, 1.667185045E9, 1.667185093E9, 1.667185141E9, 1.667185189E9, 1.667185237E9, 1.667185285E9, 1.667185333E9, 1.667185381E9, 1.667185429E9, 1.667185477E9, 1.667185525E9, 1.667185573E9, 1.667185621E9, 1.667185669E9, 1.667185717E9, 1.667185765E9, 1.667185813E9, 1.667185861E9, 1.667185909E9, 1.667185957E9, 1.667186005E9, 1.667186053E9, 1.667186101E9, 1.667186149E9, 1.66718646E9, 1.66718664E9, 1.667192466E9, 1.667192514E9, 1.667192562E9, 1.66719261E9, 1.667192658E9, 1.667192706E9, 1.667192754E9, 1.667192802E9, 1.66719285E9, 1.667192898E9, 1.667192946E9, 1.667192994E9, 1.667193042E9, 1.66719309E9, 1.667193138E9, 1.667193186E9, 1.667193234E9, 1.667193282E9, 1.66719333E9, 1.667193378E9, 1.667193426E9, 1.667193474E9, 1.667193522E9, 1.66719357E9, 1.667193618E9, 1.667193666E9, 1.667193714E9, 1.667193762E9, 1.66719381E9, 1.667193858E9, 1.667193906E9, 1.667193954E9, 1.667194002E9, 1.66719405E9, 1.667194098E9, 1.667194146E9, 1.667194194E9, 1.667194242E9, 1.66719429E9, 1.667194338E9, 1.667194386E9, 1.667194434E9, 1.667194482E9, 1.66719453E9, 1.667194578E9, 1.667194626E9, 1.667194674E9, 1.667194722E9, 1.66719477E9, 1.667194818E9, 1.667194866E9, 1.667194914E9, 1.667194962E9, 1.66719501E9, 1.667195058E9, 1.667195106E9, 1.667195154E9, 1.667195202E9, 1.66719525E9, 1.667195298E9, 1.667195346E9, 1.667195394E9, 1.667195442E9, 1.66719549E9, 1.667195538E9, 1.667195586E9, 1.667195634E9, 1.667195682E9, 1.66719573E9, 1.66719612E9, 1.6671963E9, 1.667202045E9, 1.667202093E9, 1.667202141E9, 1.667202189E9, 1.667202237E9, 1.667202285E9, 1.667202333E9, 1.667202381E9, 1.667202429E9, 1.667202477E9, 1.667202525E9, 1.667202573E9, 1.667202621E9, 1.667202669E9, 1.667202717E9, 1.667202765E9, 1.667202813E9, 1.667202861E9, 1.667202909E9, 1.667202957E9, 1.667203005E9, 1.667203053E9, 1.667203101E9, 1.667203149E9, 1.667203197E9, 1.667203245E9, 1.667203293E9, 1.667203341E9, 1.667203389E9, 1.667203437E9, 1.667203485E9, 1.667203533E9, 1.667203581E9, 1.667203629E9, 1.667203677E9, 1.667203725E9, 1.667203773E9, 1.667203821E9, 1.667203869E9, 1.667203917E9, 1.667203965E9, 1.667204013E9, 1.667204061E9, 1.667204109E9, 1.667204157E9, 1.667204205E9, 1.667204253E9, 1.667204301E9, 1.667204349E9, 1.667204397E9, 1.667204445E9, 1.667204493E9, 1.667204541E9, 1.667204589E9, 1.667204637E9, 1.667204685E9, 1.667204733E9, 1.667204781E9, 1.667204829E9, 1.667204877E9, 1.667204925E9, 1.667204973E9, 1.667205021E9, 1.667205069E9, 1.667205117E9, 1.667205165E9, 1.667205213E9, 1.667205261E9, 1.667205309E9, 1.66720566E9, 1.66720584E9, 1.667211783E9, 1.667211831E9, 1.667211879E9, 1.667211927E9, 1.667211975E9, 1.667212023E9, 1.667212071E9, 1.667212119E9, 1.667212167E9, 1.667212215E9, 1.667212263E9, 1.667212311E9, 1.667212359E9, 1.667212407E9, 1.667212455E9, 1.667212503E9, 1.667212551E9, 1.667212599E9, 1.667212647E9, 1.667212695E9, 1.667212743E9, 1.667212791E9, 1.667212839E9, 1.667212887E9, 1.667212935E9, 1.667212983E9, 1.667213031E9, 1.667213079E9, 1.667213127E9, 1.667213175E9, 1.667213223E9, 1.667213271E9, 1.667213319E9, 1.667213367E9, 1.667213415E9, 1.667213463E9, 1.667213511E9, 1.667213559E9, 1.667213607E9, 1.667213655E9, 1.667213703E9, 1.667213751E9, 1.667213799E9, 1.667213847E9, 1.667213895E9, 1.667213943E9, 1.667213991E9, 1.667214039E9, 1.667214087E9, 1.667214135E9, 1.667214183E9, 1.667214231E9, 1.667214279E9, 1.667214327E9, 1.667214375E9, 1.667214423E9, 1.667214471E9, 1.667214519E9, 1.667214567E9, 1.667214615E9, 1.667214663E9, 1.667214711E9, 1.667214759E9, 1.667214807E9, 1.667214855E9, 1.667214903E9, 1.667214951E9, 1.667214999E9, 1.66721532E9, 1.6672155E9, 1.66722127E9, 1.667221318E9, 1.667221366E9, 1.667221414E9, 1.667221462E9, 1.66722151E9, 1.667221558E9, 1.667221606E9, 1.667221654E9, 1.667221702E9, 1.66722175E9, 1.667221798E9, 1.667221846E9, 1.667221894E9, 1.667221942E9, 1.66722199E9, 1.667222038E9, 1.667222086E9, 1.667222134E9, 1.667222182E9, 1.66722223E9, 1.667222278E9, 1.667222326E9, 1.667222374E9, 1.667222422E9, 1.66722247E9, 1.667222518E9, 1.667222566E9, 1.667222614E9, 1.667222662E9, 1.66722271E9, 1.667222758E9, 1.667222806E9, 1.667222854E9, 1.667222902E9, 1.66722295E9, 1.667222998E9, 1.667223046E9, 1.667223094E9, 1.667223142E9, 1.66722319E9, 1.667223238E9, 1.667223286E9, 1.667223334E9, 1.667223382E9, 1.66722343E9, 1.667223478E9, 1.667223526E9, 1.667223574E9, 1.667223622E9, 1.66722367E9, 1.667223718E9, 1.667223766E9, 1.667223814E9, 1.667223862E9, 1.66722391E9, 1.667223958E9, 1.667224006E9, 1.667224054E9, 1.667224102E9, 1.66722415E9, 1.667224198E9, 1.667224246E9, 1.667224294E9, 1.667224342E9, 1.66722439E9, 1.667224438E9, 1.667224486E9, 1.667224534E9, 1.667224582E9, 1.66722463E9, 1.66722498E9, 1.66722516E9, 1.667231005E9, 1.667231053E9, 1.667231101E9, 1.667231149E9, 1.667231197E9, 1.667231245E9, 1.667231293E9, 1.667231341E9, 1.667231389E9, 1.667231437E9, 1.667231485E9, 1.667231533E9, 1.667231581E9, 1.667231629E9, 1.667231677E9, 1.667231725E9, 1.667231773E9, 1.667231821E9, 1.667231869E9, 1.667231917E9, 1.667231965E9, 1.667232013E9, 1.667232061E9, 1.667232109E9, 1.667232157E9, 1.667232205E9, 1.667232253E9, 1.667232301E9, 1.667232349E9, 1.667232397E9, 1.667232445E9, 1.667232493E9, 1.667232541E9, 1.667232589E9, 1.667232637E9, 1.667232685E9, 1.667232733E9, 1.667232781E9, 1.667232829E9, 1.667232877E9, 1.667232925E9, 1.667232973E9, 1.667233021E9, 1.667233069E9, 1.667233117E9, 1.667233165E9, 1.667233213E9, 1.667233261E9, 1.667233309E9, 1.667233357E9, 1.667233405E9, 1.667233453E9, 1.667233501E9, 1.667233549E9, 1.667233597E9, 1.667233645E9, 1.667233693E9, 1.667233741E9, 1.667233789E9, 1.667233837E9, 1.667233885E9, 1.667233933E9, 1.667233981E9, 1.667234029E9, 1.667234077E9, 1.667234125E9, 1.667234173E9, 1.667234221E9, 1.667234269E9, 1.667234317E9, 1.667234365E9, 1.667234413E9, 1.667234461E9, 1.667234509E9, 1.66723488E9, 1.66723506E9, 1.667240674E9, 1.667240722E9, 1.66724077E9, 1.667240818E9, 1.667240866E9, 1.667240914E9, 1.667240962E9, 1.66724101E9, 1.667241058E9, 1.667241106E9, 1.667241154E9, 1.667241202E9, 1.66724125E9, 1.667241298E9, 1.667241346E9, 1.667241394E9, 1.667241442E9, 1.66724149E9, 1.667241538E9, 1.667241586E9, 1.667241634E9, 1.667241682E9, 1.66724173E9, 1.667241778E9, 1.667241826E9, 1.667241874E9, 1.667241922E9, 1.66724197E9, 1.667242018E9, 1.667242066E9, 1.667242114E9, 1.667242162E9, 1.66724221E9, 1.667242258E9, 1.667242306E9, 1.667242354E9, 1.667242402E9, 1.66724245E9, 1.667242498E9, 1.667242546E9, 1.667242594E9, 1.667242642E9, 1.66724269E9, 1.667242738E9, 1.667242786E9, 1.667242834E9, 1.667242882E9, 1.66724293E9, 1.667242978E9, 1.667243026E9, 1.667243074E9, 1.667243122E9, 1.66724317E9, 1.667243218E9, 1.667243266E9, 1.667243314E9, 1.667243362E9, 1.66724341E9, 1.667243458E9, 1.667243506E9, 1.667243554E9, 1.667243602E9, 1.66724365E9, 1.667243698E9, 1.667243746E9, 1.667243794E9, 1.667243842E9, 1.66724389E9, 1.66724424E9, 1.66724442E9, 1.667250171E9, 1.667250219E9, 1.667250267E9, 1.667250315E9, 1.667250363E9, 1.667250411E9, 1.667250459E9, 1.667250507E9, 1.667250555E9, 1.667250603E9, 1.667250651E9, 1.667250699E9, 1.667250747E9, 1.667250795E9, 1.667250843E9, 1.667250891E9, 1.667250939E9, 1.667250987E9, 1.667251035E9, 1.667251083E9, 1.667251131E9, 1.667251179E9, 1.667251227E9, 1.667251275E9, 1.667251323E9, 1.667251371E9, 1.667251419E9, 1.667251467E9, 1.667251515E9, 1.667251563E9, 1.667251611E9, 1.667251659E9, 1.667251707E9, 1.667251755E9, 1.667251803E9, 1.667251851E9, 1.667251899E9, 1.667251947E9, 1.667251995E9, 1.667252043E9, 1.667252091E9, 1.667252139E9, 1.667252187E9, 1.667252235E9, 1.667252283E9, 1.667252331E9, 1.667252379E9, 1.667252427E9, 1.667252475E9, 1.667252523E9, 1.667252571E9, 1.667252619E9, 1.667252667E9, 1.667252715E9, 1.667252763E9, 1.667252811E9, 1.667252859E9, 1.667252907E9, 1.667252955E9, 1.667253003E9, 1.667253051E9, 1.667253099E9, 1.667253147E9, 1.667253195E9, 1.667253243E9, 1.667253291E9, 1.667253339E9, 1.6672536E9, 1.6672539E9, 1.667259686E9, 1.667259734E9, 1.667259782E9, 1.66725983E9, 1.667259878E9, 1.667259926E9, 1.667259974E9, 1.667260022E9, 1.66726007E9, 1.667260118E9, 1.667260166E9, 1.667260214E9, 1.667260262E9, 1.66726031E9, 1.667260358E9, 1.667260406E9, 1.667260454E9, 1.667260502E9, 1.66726055E9, 1.667260598E9, 1.667260646E9, 1.667260694E9, 1.667260742E9, 1.66726079E9, 1.667260838E9, 1.667260886E9, 1.667260934E9, 1.667260982E9, 1.66726103E9, 1.667261078E9, 1.667261126E9, 1.667261174E9, 1.667261222E9, 1.66726127E9, 1.667261318E9, 1.667261366E9, 1.667261414E9, 1.667261462E9, 1.66726151E9, 1.667261558E9, 1.667261606E9, 1.667261654E9, 1.667261702E9, 1.66726175E9, 1.667261798E9, 1.667261846E9, 1.667261894E9, 1.667261942E9, 1.66726199E9, 1.667262038E9, 1.667262086E9, 1.667262134E9, 1.667262182E9, 1.66726223E9, 1.667262278E9, 1.667262326E9, 1.667262374E9, 1.667262422E9, 1.66726247E9, 1.667262518E9, 1.667262566E9, 1.667262614E9, 1.667262662E9, 1.66726271E9, 1.667262758E9, 1.667262806E9, 1.667262854E9, 1.667262902E9, 1.66726295E9, 1.66726326E9, 1.66726344E9, 1.667269212E9, 1.66726926E9, 1.667269308E9, 1.667269356E9, 1.667269404E9, 1.667269452E9, 1.6672695E9, 1.667269548E9, 1.667269596E9, 1.667269644E9, 1.667269692E9, 1.66726974E9, 1.667269788E9, 1.667269836E9, 1.667269884E9, 1.667269932E9, 1.66726998E9, 1.667270028E9, 1.667270076E9, 1.667270124E9, 1.667270172E9, 1.66727022E9, 1.667270268E9, 1.667270316E9, 1.667270364E9, 1.667270412E9, 1.66727046E9, 1.667270508E9, 1.667270556E9, 1.667270604E9, 1.667270652E9, 1.6672707E9, 1.667270748E9, 1.667270796E9, 1.667270844E9, 1.667270892E9, 1.66727094E9, 1.667270988E9, 1.667271036E9, 1.667271084E9, 1.667271132E9, 1.66727118E9, 1.667271228E9, 1.667271276E9, 1.667271324E9, 1.667271372E9, 1.66727142E9, 1.667271468E9, 1.667271516E9, 1.667271564E9, 1.667271612E9, 1.66727166E9, 1.667271708E9, 1.667271756E9, 1.667271804E9, 1.667271852E9, 1.6672719E9, 1.667271948E9, 1.667271996E9, 1.667272044E9, 1.667272092E9, 1.66727214E9, 1.667272188E9, 1.667272236E9, 1.667272284E9, 1.667272332E9, 1.66727238E9, 1.667272428E9, 1.667272476E9, 1.667272524E9, 1.667272572E9, 1.66727262E9, 1.66727292E9, 1.6672731E9, 1.667278872E9, 1.66727892E9, 1.667278968E9, 1.667279016E9, 1.667279064E9, 1.667279112E9, 1.66727916E9, 1.667279208E9, 1.667279256E9, 1.667279304E9, 1.667279352E9, 1.6672794E9, 1.667279448E9, 1.667279496E9, 1.667279544E9, 1.667279592E9, 1.66727964E9, 1.667279688E9, 1.667279736E9, 1.667279784E9, 1.667279832E9, 1.66727988E9, 1.667279928E9, 1.667279976E9, 1.667280024E9, 1.667280072E9, 1.66728012E9, 1.667280168E9, 1.667280216E9, 1.667280264E9, 1.667280312E9, 1.66728036E9, 1.667280408E9, 1.667280456E9, 1.667280504E9, 1.667280552E9, 1.6672806E9, 1.667280648E9, 1.667280696E9, 1.667280744E9, 1.667280792E9, 1.66728084E9, 1.667280888E9, 1.667280936E9, 1.667280984E9, 1.667281032E9, 1.66728108E9, 1.667281128E9, 1.667281176E9, 1.667281224E9, 1.667281272E9, 1.66728132E9, 1.667281368E9, 1.667281416E9, 1.667281464E9, 1.667281512E9, 1.66728156E9, 1.667281608E9, 1.667281656E9, 1.667281704E9, 1.667281752E9, 1.6672818E9, 1.667281848E9, 1.667281896E9, 1.667281944E9, 1.667281992E9, 1.66728204E9, 1.66728234E9, 1.66728252E9, 1.667288574E9, 1.667288622E9, 1.66728867E9, 1.667288718E9, 1.667288766E9, 1.667288814E9, 1.667288862E9, 1.66728891E9, 1.667288958E9, 1.667289006E9, 1.667289054E9, 1.667289102E9, 1.66728915E9, 1.667289198E9, 1.667289246E9, 1.667289294E9, 1.667289342E9, 1.66728939E9, 1.667289438E9, 1.667289486E9, 1.667289534E9, 1.667289582E9, 1.66728963E9, 1.667289678E9, 1.667289726E9, 1.667289774E9, 1.667289822E9, 1.66728987E9, 1.667289918E9, 1.667289966E9, 1.667290014E9, 1.667290062E9, 1.66729011E9, 1.667290158E9, 1.667290206E9, 1.667290254E9, 1.667290302E9, 1.66729035E9, 1.667290398E9, 1.667290446E9, 1.667290494E9, 1.667290542E9, 1.66729059E9, 1.667290638E9, 1.667290686E9, 1.667290734E9, 1.667290782E9, 1.66729083E9, 1.667290878E9, 1.667290926E9, 1.667290974E9, 1.667291022E9, 1.66729107E9, 1.667291118E9, 1.667291166E9, 1.667291214E9, 1.667291262E9, 1.66729131E9, 1.667291358E9, 1.667291406E9, 1.667291454E9, 1.667291502E9, 1.66729155E9, 1.667291598E9, 1.667291646E9, 1.667291694E9, 1.667291742E9, 1.66729179E9, 1.66729212E9, 1.6672923E9, 1.667298051E9, 1.667298099E9, 1.667298147E9, 1.667298195E9, 1.667298243E9, 1.667298291E9, 1.667298339E9, 1.667298387E9, 1.667298435E9, 1.667298483E9, 1.667298531E9, 1.667298579E9, 1.667298627E9, 1.667298675E9, 1.667298723E9, 1.667298771E9, 1.667298819E9, 1.667298867E9, 1.667298915E9, 1.667298963E9, 1.667299011E9, 1.667299059E9, 1.667299107E9, 1.667299155E9, 1.667299203E9, 1.667299251E9, 1.667299299E9, 1.667299347E9, 1.667299395E9, 1.667299443E9, 1.667299491E9, 1.667299539E9, 1.667299587E9, 1.667299635E9, 1.667299683E9, 1.667299731E9, 1.667299779E9, 1.667299827E9, 1.667299875E9, 1.667299923E9, 1.667299971E9, 1.667300019E9, 1.667300067E9, 1.667300115E9, 1.667300163E9, 1.667300211E9, 1.667300259E9, 1.667300307E9, 1.667300355E9, 1.667300403E9, 1.667300451E9, 1.667300499E9, 1.667300547E9, 1.667300595E9, 1.667300643E9, 1.667300691E9, 1.667300739E9, 1.667300787E9, 1.667300835E9, 1.667300883E9, 1.667300931E9, 1.667300979E9, 1.667301027E9, 1.667301075E9, 1.667301123E9, 1.667301171E9, 1.667301219E9, 1.66730148E9, 1.66730172E9, 1.667307537E9, 1.667307585E9, 1.667307633E9, 1.667307681E9, 1.667307729E9, 1.667307777E9, 1.667307825E9, 1.667307873E9, 1.667307921E9, 1.667307969E9, 1.667308017E9, 1.667308065E9, 1.667308113E9, 1.667308161E9, 1.667308209E9, 1.667308257E9, 1.667308305E9, 1.667308353E9, 1.667308401E9, 1.667308449E9, 1.667308497E9, 1.667308545E9, 1.667308593E9, 1.667308641E9, 1.667308689E9, 1.667308737E9, 1.667308785E9, 1.667308833E9, 1.667308881E9, 1.667308929E9, 1.667308977E9, 1.667309025E9, 1.667309073E9, 1.667309121E9, 1.667309169E9, 1.667309217E9, 1.667309265E9, 1.667309313E9, 1.667309361E9, 1.667309409E9, 1.667309457E9, 1.667309505E9, 1.667309553E9, 1.667309601E9, 1.667309649E9, 1.667309697E9, 1.667309745E9, 1.667309793E9, 1.667309841E9, 1.667309889E9, 1.667309937E9, 1.667309985E9, 1.667310033E9, 1.667310081E9, 1.667310129E9, 1.667310177E9, 1.667310225E9, 1.667310273E9, 1.667310321E9, 1.667310369E9, 1.667310417E9, 1.667310465E9, 1.667310513E9, 1.667310561E9, 1.667310609E9, 1.667310657E9, 1.667310705E9, 1.667310753E9, 1.667310801E9, 1.667310849E9, 1.66731114E9, 1.66731132E9, 1.667317123E9, 1.667317171E9, 1.667317219E9, 1.667317267E9, 1.667317315E9, 1.667317363E9, 1.667317411E9, 1.667317459E9, 1.667317507E9, 1.667317555E9, 1.667317603E9, 1.667317651E9, 1.667317699E9, 1.667317747E9, 1.667317795E9, 1.667317843E9, 1.667317891E9, 1.667317939E9, 1.667317987E9, 1.667318035E9, 1.667318083E9, 1.667318131E9, 1.667318179E9, 1.667318227E9, 1.667318275E9, 1.667318323E9, 1.667318371E9, 1.667318419E9, 1.667318467E9, 1.667318515E9, 1.667318563E9, 1.667318611E9, 1.667318659E9, 1.667318707E9, 1.667318755E9, 1.667318803E9, 1.667318851E9, 1.667318899E9, 1.667318947E9, 1.667318995E9, 1.667319043E9, 1.667319091E9, 1.667319139E9, 1.667319187E9, 1.667319235E9, 1.667319283E9, 1.667319331E9, 1.667319379E9, 1.667319427E9, 1.667319475E9, 1.667319523E9, 1.667319571E9, 1.667319619E9, 1.667319667E9, 1.667319715E9, 1.667319763E9, 1.667319811E9, 1.667319859E9, 1.667319907E9, 1.667319955E9, 1.667320003E9, 1.667320051E9, 1.667320099E9, 1.667320147E9, 1.667320195E9, 1.667320243E9, 1.667320291E9, 1.667320339E9, 1.66732074E9, 1.66732092E9, 1.667326561E9, 1.667326609E9, 1.667326657E9, 1.667326705E9, 1.667326753E9, 1.667326801E9, 1.667326849E9, 1.667326897E9, 1.667326945E9, 1.667326993E9, 1.667327041E9, 1.667327089E9, 1.667327137E9, 1.667327185E9, 1.667327233E9, 1.667327281E9, 1.667327329E9, 1.667327377E9, 1.667327425E9, 1.667327473E9, 1.667327521E9, 1.667327569E9, 1.667327617E9, 1.667327665E9, 1.667327713E9, 1.667327761E9, 1.667327809E9, 1.667327857E9, 1.667327905E9, 1.667327953E9, 1.667328001E9, 1.667328049E9, 1.667328097E9, 1.667328145E9, 1.667328193E9, 1.667328241E9, 1.667328289E9, 1.667328337E9, 1.667328385E9, 1.667328433E9, 1.667328481E9, 1.667328529E9, 1.667328577E9, 1.667328625E9, 1.667328673E9, 1.667328721E9, 1.667328769E9, 1.667328817E9, 1.667328865E9, 1.667328913E9, 1.667328961E9, 1.667329009E9, 1.667329057E9, 1.667329105E9, 1.667329153E9, 1.667329201E9, 1.667329249E9, 1.667329297E9, 1.667329345E9, 1.667329393E9, 1.667329441E9, 1.667329489E9, 1.667329537E9, 1.667329585E9, 1.667329633E9, 1.667329681E9, 1.667329729E9, 1.66733004E9, 1.66733022E9, 1.667335772E9, 1.66733582E9, 1.667335868E9, 1.667335916E9, 1.667335964E9, 1.667336012E9, 1.66733606E9, 1.667336108E9, 1.667336156E9, 1.667336204E9, 1.667336252E9, 1.6673363E9, 1.667336348E9, 1.667336396E9, 1.667336444E9, 1.667336492E9, 1.66733654E9, 1.667336588E9, 1.667336636E9, 1.667336684E9, 1.667336732E9, 1.66733678E9, 1.667336828E9, 1.667336876E9, 1.667336924E9, 1.667336972E9, 1.66733702E9, 1.667337068E9, 1.667337116E9, 1.667337164E9, 1.667337212E9, 1.66733726E9, 1.667337308E9, 1.667337356E9, 1.667337404E9, 1.667337452E9, 1.6673375E9, 1.667337548E9, 1.667337596E9, 1.667337644E9, 1.667337692E9, 1.66733774E9, 1.667337788E9, 1.667337836E9, 1.667337884E9, 1.667337932E9, 1.66733798E9, 1.667338028E9, 1.667338076E9, 1.667338124E9, 1.667338172E9, 1.66733822E9, 1.667338268E9, 1.667338316E9, 1.667338364E9, 1.667338412E9, 1.66733846E9, 1.667338508E9, 1.667338556E9, 1.667338604E9, 1.667338652E9, 1.6673387E9, 1.667338748E9, 1.667338796E9, 1.667338844E9, 1.667338892E9, 1.66733894E9, 1.667338988E9, 1.667339036E9, 1.667339084E9, 1.667339132E9, 1.66733918E9, 1.66733958E9, 1.66733976E9, 1.667345516E9, 1.667345564E9, 1.667345612E9, 1.66734566E9, 1.667345708E9, 1.667345756E9, 1.667345804E9, 1.667345852E9, 1.6673459E9, 1.667345948E9, 1.667345996E9, 1.667346044E9, 1.667346092E9, 1.66734614E9, 1.667346188E9, 1.667346236E9, 1.667346284E9, 1.667346332E9, 1.66734638E9, 1.667346428E9, 1.667346476E9, 1.667346524E9, 1.667346572E9, 1.66734662E9, 1.667346668E9, 1.667346716E9, 1.667346764E9, 1.667346812E9, 1.66734686E9, 1.667346908E9, 1.667346956E9, 1.667347004E9, 1.667347052E9, 1.6673471E9, 1.667347148E9, 1.667347196E9, 1.667347244E9, 1.667347292E9, 1.66734734E9, 1.667347388E9, 1.667347436E9, 1.667347484E9, 1.667347532E9, 1.66734758E9, 1.667347628E9, 1.667347676E9, 1.667347724E9, 1.667347772E9, 1.66734782E9, 1.667347868E9, 1.667347916E9, 1.667347964E9, 1.667348012E9, 1.66734806E9, 1.667348108E9, 1.667348156E9, 1.667348204E9, 1.667348252E9, 1.6673483E9, 1.667348348E9, 1.667348396E9, 1.667348444E9, 1.667348492E9, 1.66734854E9, 1.667348588E9, 1.667348636E9, 1.667348684E9, 1.667348732E9, 1.66734878E9, 1.66734918E9, 1.667349181E9, 1.667354913E9, 1.667354961E9, 1.667355009E9, 1.667355057E9, 1.667355105E9, 1.667355153E9, 1.667355201E9, 1.667355249E9, 1.667355297E9, 1.667355345E9, 1.667355393E9, 1.667355441E9, 1.667355489E9, 1.667355537E9, 1.667355585E9, 1.667355633E9, 1.667355681E9, 1.667355729E9, 1.667355777E9, 1.667355825E9, 1.667355873E9, 1.667355921E9, 1.667355969E9, 1.667356017E9, 1.667356065E9, 1.667356113E9, 1.667356161E9, 1.667356209E9, 1.667356257E9, 1.667356305E9, 1.667356353E9, 1.667356401E9, 1.667356449E9, 1.667356497E9, 1.667356545E9, 1.667356593E9, 1.667356641E9, 1.667356689E9, 1.667356737E9, 1.667356785E9, 1.667356833E9, 1.667356881E9, 1.667356929E9, 1.667356977E9, 1.667357025E9, 1.667357073E9, 1.667357121E9, 1.667357169E9, 1.667357217E9, 1.667357265E9, 1.667357313E9, 1.667357361E9, 1.667357409E9, 1.667357457E9, 1.667357505E9, 1.667357553E9, 1.667357601E9, 1.667357649E9, 1.667357697E9, 1.667357745E9, 1.667357793E9, 1.667357841E9, 1.667357889E9, 1.667357937E9, 1.667357985E9, 1.667358033E9, 1.667358081E9, 1.667358129E9, 1.66735842E9, 1.6673586E9, 1.667364289E9, 1.667364337E9, 1.667364385E9, 1.667364433E9, 1.667364481E9, 1.667364529E9, 1.667364577E9, 1.667364625E9, 1.667364673E9, 1.667364721E9, 1.667364769E9, 1.667364817E9, 1.667364865E9, 1.667364913E9, 1.667364961E9, 1.667365009E9, 1.667365057E9, 1.667365105E9, 1.667365153E9, 1.667365201E9, 1.667365249E9, 1.667365297E9, 1.667365345E9, 1.667365393E9, 1.667365441E9, 1.667365489E9, 1.667365537E9, 1.667365585E9, 1.667365633E9, 1.667365681E9, 1.667365729E9, 1.667365777E9, 1.667365825E9, 1.667365873E9, 1.667365921E9, 1.667365969E9, 1.667366017E9, 1.667366065E9, 1.667366113E9, 1.667366161E9, 1.667366209E9, 1.667366257E9, 1.667366305E9, 1.667366353E9, 1.667366401E9, 1.667366449E9, 1.667366497E9, 1.667366545E9, 1.667366593E9, 1.667366641E9, 1.667366689E9, 1.667366737E9, 1.667366785E9, 1.667366833E9, 1.667366881E9, 1.667366929E9, 1.667366977E9, 1.667367025E9, 1.667367073E9, 1.667367121E9, 1.667367169E9, 1.667367217E9, 1.667367265E9, 1.667367313E9, 1.667367361E9, 1.667367409E9, 1.667367457E9, 1.667367505E9, 1.667367553E9, 1.667367601E9, 1.667367649E9, 1.66736796E9, 1.66736814E9, 1.667373703E9, 1.667373751E9, 1.667373799E9, 1.667373847E9, 1.667373895E9, 1.667373943E9, 1.667373991E9, 1.667374039E9, 1.667374087E9, 1.667374135E9, 1.667374183E9, 1.667374231E9, 1.667374279E9, 1.667374327E9, 1.667374375E9, 1.667374423E9, 1.667374471E9, 1.667374519E9, 1.667374567E9, 1.667374615E9, 1.667374663E9, 1.667374711E9, 1.667374759E9, 1.667374807E9, 1.667374855E9, 1.667374903E9, 1.667374951E9, 1.667374999E9, 1.667375047E9, 1.667375095E9, 1.667375143E9, 1.667375191E9, 1.667375239E9, 1.667375287E9, 1.667375335E9, 1.667375383E9, 1.667375431E9, 1.667375479E9, 1.667375527E9, 1.667375575E9, 1.667375623E9, 1.667375671E9, 1.667375719E9, 1.667375767E9, 1.667375815E9, 1.667375863E9, 1.667375911E9, 1.667375959E9, 1.667376007E9, 1.667376055E9, 1.667376103E9, 1.667376151E9, 1.667376199E9, 1.667376247E9, 1.667376295E9, 1.667376343E9, 1.667376391E9, 1.667376439E9, 1.667376487E9, 1.667376535E9, 1.667376583E9, 1.667376631E9, 1.667376679E9, 1.667376727E9, 1.667376775E9, 1.667376823E9, 1.667376871E9, 1.667376919E9, 1.66737732E9, 1.6673775E9, 1.667383184E9, 1.667383232E9, 1.66738328E9, 1.667383328E9, 1.667383376E9, 1.667383424E9, 1.667383472E9, 1.66738352E9, 1.667383568E9, 1.667383616E9, 1.667383664E9, 1.667383712E9, 1.66738376E9, 1.667383808E9, 1.667383856E9, 1.667383904E9, 1.667383952E9, 1.667384E9, 1.667384048E9, 1.667384096E9, 1.667384144E9, 1.667384192E9, 1.66738424E9, 1.667384288E9, 1.667384336E9, 1.667384384E9, 1.667384432E9, 1.66738448E9, 1.667384528E9, 1.667384576E9, 1.667384624E9, 1.667384672E9, 1.66738472E9, 1.667384768E9, 1.667384816E9, 1.667384864E9, 1.667384912E9, 1.66738496E9, 1.667385008E9, 1.667385056E9, 1.667385104E9, 1.667385152E9, 1.6673852E9, 1.667385248E9, 1.667385296E9, 1.667385344E9, 1.667385392E9, 1.66738544E9, 1.667385488E9, 1.667385536E9, 1.667385584E9, 1.667385632E9, 1.66738568E9, 1.667385728E9, 1.667385776E9, 1.667385824E9, 1.667385872E9, 1.66738592E9, 1.667385968E9, 1.667386016E9, 1.667386064E9, 1.667386112E9, 1.66738616E9, 1.667386208E9, 1.667386256E9, 1.667386304E9, 1.667386352E9, 1.6673864E9, 1.66738668E9, 1.66738686E9, 1.667392473E9, 1.667392521E9, 1.667392569E9, 1.667392617E9, 1.667392665E9, 1.667392713E9, 1.667392761E9, 1.667392809E9, 1.667392857E9, 1.667392905E9, 1.667392953E9, 1.667393001E9, 1.667393049E9, 1.667393097E9, 1.667393145E9, 1.667393193E9, 1.667393241E9, 1.667393289E9, 1.667393337E9, 1.667393385E9, 1.667393433E9, 1.667393481E9, 1.667393529E9, 1.667393577E9, 1.667393625E9, 1.667393673E9, 1.667393721E9, 1.667393769E9, 1.667393817E9, 1.667393865E9, 1.667393913E9, 1.667393961E9, 1.667394009E9, 1.667394057E9, 1.667394105E9, 1.667394153E9, 1.667394201E9, 1.667394249E9, 1.667394297E9, 1.667394345E9, 1.667394393E9, 1.667394441E9, 1.667394489E9, 1.667394537E9, 1.667394585E9, 1.667394633E9, 1.667394681E9, 1.667394729E9, 1.667394777E9, 1.667394825E9, 1.667394873E9, 1.667394921E9, 1.667394969E9, 1.667395017E9, 1.667395065E9, 1.667395113E9, 1.667395161E9, 1.667395209E9, 1.667395257E9, 1.667395305E9, 1.667395353E9, 1.667395401E9, 1.667395449E9, 1.667395497E9, 1.667395545E9, 1.667395593E9, 1.667395641E9, 1.667395689E9, 1.667395737E9, 1.667395785E9, 1.667395833E9, 1.667395881E9, 1.667395929E9, 1.66739616E9, 1.66739634E9, 1.6674024E9, 1.667402448E9, 1.667402496E9, 1.667402544E9, 1.667402592E9, 1.66740264E9, 1.667402688E9, 1.667402736E9, 1.667402784E9, 1.667402832E9, 1.66740288E9, 1.667402928E9, 1.667402976E9, 1.667403024E9, 1.667403072E9, 1.66740312E9, 1.667403168E9, 1.667403216E9, 1.667403264E9, 1.667403312E9, 1.66740336E9, 1.667403408E9, 1.667403456E9, 1.667403504E9, 1.667403552E9, 1.6674036E9, 1.667403648E9, 1.667403696E9, 1.667403744E9, 1.667403792E9, 1.66740384E9, 1.667403888E9, 1.667403936E9, 1.667403984E9, 1.667404032E9, 1.66740408E9, 1.667404128E9, 1.667404176E9, 1.667404224E9, 1.667404272E9, 1.66740432E9, 1.667404368E9, 1.667404416E9, 1.667404464E9, 1.667404512E9, 1.66740456E9, 1.667404608E9, 1.667404656E9, 1.667404704E9, 1.667404752E9, 1.6674048E9, 1.667404848E9, 1.667404896E9, 1.667404944E9, 1.667404992E9, 1.66740504E9, 1.667405088E9, 1.667405136E9, 1.667405184E9, 1.667405232E9, 1.66740528E9, 1.667405328E9, 1.667405376E9, 1.667405424E9, 1.667405472E9, 1.66740552E9, 1.66740588E9, 1.667405881E9, 1.667411575E9, 1.667411623E9, 1.667411671E9, 1.667411719E9, 1.667411767E9, 1.667411815E9, 1.667411863E9, 1.667411911E9, 1.667411959E9, 1.667412007E9, 1.667412055E9, 1.667412103E9, 1.667412151E9, 1.667412199E9, 1.667412247E9, 1.667412295E9, 1.667412343E9, 1.667412391E9, 1.667412439E9, 1.667412487E9, 1.667412535E9, 1.667412583E9, 1.667412631E9, 1.667412679E9, 1.667412727E9, 1.667412775E9, 1.667412823E9, 1.667412871E9, 1.667412919E9, 1.667412967E9, 1.667413015E9, 1.667413063E9, 1.667413111E9, 1.667413159E9, 1.667413207E9, 1.667413255E9, 1.667413303E9, 1.667413351E9, 1.667413399E9, 1.667413447E9, 1.667413495E9, 1.667413543E9, 1.667413591E9, 1.667413639E9, 1.667413687E9, 1.667413735E9, 1.667413783E9, 1.667413831E9, 1.667413879E9, 1.667413927E9, 1.667413975E9, 1.667414023E9, 1.667414071E9, 1.667414119E9, 1.667414167E9, 1.667414215E9, 1.667414263E9, 1.667414311E9, 1.667414359E9, 1.667414407E9, 1.667414455E9, 1.667414503E9, 1.667414551E9, 1.667414599E9, 1.667414647E9, 1.667414695E9, 1.667414743E9, 1.667414791E9, 1.667414839E9, 1.66741512E9, 1.6674153E9, 1.667420981E9, 1.667421029E9, 1.667421077E9, 1.667421125E9, 1.667421173E9, 1.667421221E9, 1.667421269E9, 1.667421317E9, 1.667421365E9, 1.667421413E9, 1.667421461E9, 1.667421509E9, 1.667421557E9, 1.667421605E9, 1.667421653E9, 1.667421701E9, 1.667421749E9, 1.667421797E9, 1.667421845E9, 1.667421893E9, 1.667421941E9, 1.667421989E9, 1.667422037E9, 1.667422085E9, 1.667422133E9, 1.667422181E9, 1.667422229E9, 1.667422277E9, 1.667422325E9, 1.667422373E9, 1.667422421E9, 1.667422469E9, 1.667422517E9, 1.667422565E9, 1.667422613E9, 1.667422661E9, 1.667422709E9, 1.667422757E9, 1.667422805E9, 1.667422853E9, 1.667422901E9, 1.667422949E9, 1.667422997E9, 1.667423045E9, 1.667423093E9, 1.667423141E9, 1.667423189E9, 1.667423237E9, 1.667423285E9, 1.667423333E9, 1.667423381E9, 1.667423429E9, 1.667423477E9, 1.667423525E9, 1.667423573E9, 1.667423621E9, 1.667423669E9, 1.667423717E9, 1.667423765E9, 1.667423813E9, 1.667423861E9, 1.667423909E9, 1.667423957E9, 1.667424005E9, 1.667424053E9, 1.667424101E9, 1.667424149E9, 1.667424197E9, 1.667424245E9, 1.667424293E9, 1.667424341E9, 1.667424389E9, 1.66742472E9, 1.6674249E9, 1.667430619E9, 1.667430667E9, 1.667430715E9, 1.667430763E9, 1.667430811E9, 1.667430859E9, 1.667430907E9, 1.667430955E9, 1.667431003E9, 1.667431051E9, 1.667431099E9, 1.667431147E9, 1.667431195E9, 1.667431243E9, 1.667431291E9, 1.667431339E9, 1.667431387E9, 1.667431435E9, 1.667431483E9, 1.667431531E9, 1.667431579E9, 1.667431627E9, 1.667431675E9, 1.667431723E9, 1.667431771E9, 1.667431819E9, 1.667431867E9, 1.667431915E9, 1.667431963E9, 1.667432011E9, 1.667432059E9, 1.667432107E9, 1.667432155E9, 1.667432203E9, 1.667432251E9, 1.667432299E9, 1.667432347E9, 1.667432395E9, 1.667432443E9, 1.667432491E9, 1.667432539E9, 1.667432587E9, 1.667432635E9, 1.667432683E9, 1.667432731E9, 1.667432779E9, 1.667432827E9, 1.667432875E9, 1.667432923E9, 1.667432971E9, 1.667433019E9, 1.667433067E9, 1.667433115E9, 1.667433163E9, 1.667433211E9, 1.667433259E9, 1.667433307E9, 1.667433355E9, 1.667433403E9, 1.667433451E9, 1.667433499E9, 1.667433547E9, 1.667433595E9, 1.667433643E9, 1.667433691E9, 1.667433739E9, 1.667433787E9, 1.667433835E9, 1.667433883E9, 1.667433931E9, 1.667433979E9, 1.66743432E9, 1.6674345E9, 1.667440053E9, 1.667440101E9, 1.667440149E9, 1.667440197E9, 1.667440245E9, 1.667440293E9, 1.667440341E9, 1.667440389E9, 1.667440437E9, 1.667440485E9, 1.667440533E9, 1.667440581E9, 1.667440629E9, 1.667440677E9, 1.667440725E9, 1.667440773E9, 1.667440821E9, 1.667440869E9, 1.667440917E9, 1.667440965E9, 1.667441013E9, 1.667441061E9, 1.667441109E9, 1.667441157E9, 1.667441205E9, 1.667441253E9, 1.667441301E9, 1.667441349E9, 1.667441397E9, 1.667441445E9, 1.667441493E9, 1.667441541E9, 1.667441589E9, 1.667441637E9, 1.667441685E9, 1.667441733E9, 1.667441781E9, 1.667441829E9, 1.667441877E9, 1.667441925E9, 1.667441973E9, 1.667442021E9, 1.667442069E9, 1.667442117E9, 1.667442165E9, 1.667442213E9, 1.667442261E9, 1.667442309E9, 1.667442357E9, 1.667442405E9, 1.667442453E9, 1.667442501E9, 1.667442549E9, 1.667442597E9, 1.667442645E9, 1.667442693E9, 1.667442741E9, 1.667442789E9, 1.667442837E9, 1.667442885E9, 1.667442933E9, 1.667442981E9, 1.667443029E9, 1.667443077E9, 1.667443125E9, 1.667443173E9, 1.667443221E9, 1.667443269E9, 1.667443317E9, 1.667443365E9, 1.667443413E9, 1.667443461E9, 1.667443509E9, 1.66744374E9, 1.66744392E9, 1.667449653E9, 1.667449701E9, 1.667449749E9, 1.667449797E9, 1.667449845E9, 1.667449893E9, 1.667449941E9, 1.667449989E9, 1.667450037E9, 1.667450085E9, 1.667450133E9, 1.667450181E9, 1.667450229E9, 1.667450277E9, 1.667450325E9, 1.667450373E9, 1.667450421E9, 1.667450469E9, 1.667450517E9, 1.667450565E9, 1.667450613E9, 1.667450661E9, 1.667450709E9, 1.667450757E9, 1.667450805E9, 1.667450853E9, 1.667450901E9, 1.667450949E9, 1.667450997E9, 1.667451045E9, 1.667451093E9, 1.667451141E9, 1.667451189E9, 1.667451237E9, 1.667451285E9, 1.667451333E9, 1.667451381E9, 1.667451429E9, 1.667451477E9, 1.667451525E9, 1.667451573E9, 1.667451621E9, 1.667451669E9, 1.667451717E9, 1.667451765E9, 1.667451813E9, 1.667451861E9, 1.667451909E9, 1.667451957E9, 1.667452005E9, 1.667452053E9, 1.667452101E9, 1.667452149E9, 1.667452197E9, 1.667452245E9, 1.667452293E9, 1.667452341E9, 1.667452389E9, 1.667452437E9, 1.667452485E9, 1.667452533E9, 1.667452581E9, 1.667452629E9, 1.667452677E9, 1.667452725E9, 1.667452773E9, 1.667452821E9, 1.667452869E9, 1.667452917E9, 1.667452965E9, 1.667453013E9, 1.667453061E9, 1.667453109E9, 1.6674534E9, 1.66745358E9, 1.667459184E9, 1.667459232E9, 1.66745928E9, 1.667459328E9, 1.667459376E9, 1.667459424E9, 1.667459472E9, 1.66745952E9, 1.667459568E9, 1.667459616E9, 1.667459664E9, 1.667459712E9, 1.66745976E9, 1.667459808E9, 1.667459856E9, 1.667459904E9, 1.667459952E9, 1.66746E9, 1.667460048E9, 1.667460096E9, 1.667460144E9, 1.667460192E9, 1.66746024E9, 1.667460288E9, 1.667460336E9, 1.667460384E9, 1.667460432E9, 1.66746048E9, 1.667460528E9, 1.667460576E9, 1.667460624E9, 1.667460672E9, 1.66746072E9, 1.667460768E9, 1.667460816E9, 1.667460864E9, 1.667460912E9, 1.66746096E9, 1.667461008E9, 1.667461056E9, 1.667461104E9, 1.667461152E9, 1.6674612E9, 1.667461248E9, 1.667461296E9, 1.667461344E9, 1.667461392E9, 1.66746144E9, 1.667461488E9, 1.667461536E9, 1.667461584E9, 1.667461632E9, 1.66746168E9, 1.667461728E9, 1.667461776E9, 1.667461824E9, 1.667461872E9, 1.66746192E9, 1.667461968E9, 1.667462016E9, 1.667462064E9, 1.667462112E9, 1.66746216E9, 1.667462208E9, 1.667462256E9, 1.667462304E9, 1.667462352E9, 1.6674624E9, 1.66746276E9, 1.66746294E9, 1.667468544E9, 1.667468592E9, 1.66746864E9, 1.667468688E9, 1.667468736E9, 1.667468784E9, 1.667468832E9, 1.66746888E9, 1.667468928E9, 1.667468976E9, 1.667469024E9, 1.667469072E9, 1.66746912E9, 1.667469168E9, 1.667469216E9, 1.667469264E9, 1.667469312E9, 1.66746936E9, 1.667469408E9, 1.667469456E9, 1.667469504E9, 1.667469552E9, 1.6674696E9, 1.667469648E9, 1.667469696E9, 1.667469744E9, 1.667469792E9, 1.66746984E9, 1.667469888E9, 1.667469936E9, 1.667469984E9, 1.667470032E9, 1.66747008E9, 1.667470128E9, 1.667470176E9, 1.667470224E9, 1.667470272E9, 1.66747032E9, 1.667470368E9, 1.667470416E9, 1.667470464E9, 1.667470512E9, 1.66747056E9, 1.667470608E9, 1.667470656E9, 1.667470704E9, 1.667470752E9, 1.6674708E9, 1.667470848E9, 1.667470896E9, 1.667470944E9, 1.667470992E9, 1.66747104E9, 1.667471088E9, 1.667471136E9, 1.667471184E9, 1.667471232E9, 1.66747128E9, 1.667471328E9, 1.667471376E9, 1.667471424E9, 1.667471472E9, 1.66747152E9, 1.667471568E9, 1.667471616E9, 1.667471664E9, 1.667471712E9, 1.66747176E9, 1.66747206E9, 1.66747224E9, 1.667477954E9, 1.667478002E9, 1.66747805E9, 1.667478098E9, 1.667478146E9, 1.667478194E9, 1.667478242E9, 1.66747829E9, 1.667478338E9, 1.667478386E9, 1.667478434E9, 1.667478482E9, 1.66747853E9, 1.667478578E9, 1.667478626E9, 1.667478674E9, 1.667478722E9, 1.66747877E9, 1.667478818E9, 1.667478866E9, 1.667478914E9, 1.667478962E9, 1.66747901E9, 1.667479058E9, 1.667479106E9, 1.667479154E9, 1.667479202E9, 1.66747925E9, 1.667479298E9, 1.667479346E9, 1.667479394E9, 1.667479442E9, 1.66747949E9, 1.667479538E9, 1.667479586E9, 1.667479634E9, 1.667479682E9, 1.66747973E9, 1.667479778E9, 1.667479826E9, 1.667479874E9, 1.667479922E9, 1.66747997E9, 1.667480018E9, 1.667480066E9, 1.667480114E9, 1.667480162E9, 1.66748021E9, 1.667480258E9, 1.667480306E9, 1.667480354E9, 1.667480402E9, 1.66748045E9, 1.667480498E9, 1.667480546E9, 1.667480594E9, 1.667480642E9, 1.66748069E9, 1.667480738E9, 1.667480786E9, 1.667480834E9, 1.667480882E9, 1.66748093E9, 1.667480978E9, 1.667481026E9, 1.667481074E9, 1.667481122E9, 1.66748117E9, 1.66748148E9, 1.66748166E9, 1.667487566E9, 1.667487614E9, 1.667487662E9, 1.66748771E9, 1.667487758E9, 1.667487806E9, 1.667487854E9, 1.667487902E9, 1.66748795E9, 1.667487998E9, 1.667488046E9, 1.667488094E9, 1.667488142E9, 1.66748819E9, 1.667488238E9, 1.667488286E9, 1.667488334E9, 1.667488382E9, 1.66748843E9, 1.667488478E9, 1.667488526E9, 1.667488574E9, 1.667488622E9, 1.66748867E9, 1.667488718E9, 1.667488766E9, 1.667488814E9, 1.667488862E9, 1.66748891E9, 1.667488958E9, 1.667489006E9, 1.667489054E9, 1.667489102E9, 1.66748915E9, 1.667489198E9, 1.667489246E9, 1.667489294E9, 1.667489342E9, 1.66748939E9, 1.667489438E9, 1.667489486E9, 1.667489534E9, 1.667489582E9, 1.66748963E9, 1.667489678E9, 1.667489726E9, 1.667489774E9, 1.667489822E9, 1.66748987E9, 1.667489918E9, 1.667489966E9, 1.667490014E9, 1.667490062E9, 1.66749011E9, 1.667490158E9, 1.667490206E9, 1.667490254E9, 1.667490302E9, 1.66749035E9, 1.667490398E9, 1.667490446E9, 1.667490494E9, 1.667490542E9, 1.66749059E9, 1.667490638E9, 1.667490686E9, 1.667490734E9, 1.667490782E9, 1.66749083E9, 1.66749114E9, 1.66749132E9, 1.66749688E9, 1.667496928E9, 1.667496976E9, 1.667497024E9, 1.667497072E9, 1.66749712E9, 1.667497168E9, 1.667497216E9, 1.667497264E9, 1.667497312E9, 1.66749736E9, 1.667497408E9, 1.667497456E9, 1.667497504E9, 1.667497552E9, 1.6674976E9, 1.667497648E9, 1.667497696E9, 1.667497744E9, 1.667497792E9, 1.66749784E9, 1.667497888E9, 1.667497936E9, 1.667497984E9, 1.667498032E9, 1.66749808E9, 1.667498128E9, 1.667498176E9, 1.667498224E9, 1.667498272E9, 1.66749832E9, 1.667498368E9, 1.667498416E9, 1.667498464E9, 1.667498512E9, 1.66749856E9, 1.667498608E9, 1.667498656E9, 1.667498704E9, 1.667498752E9, 1.6674988E9, 1.667498848E9, 1.667498896E9, 1.667498944E9, 1.667498992E9, 1.66749904E9, 1.667499088E9, 1.667499136E9, 1.667499184E9, 1.667499232E9, 1.66749928E9, 1.667499328E9, 1.667499376E9, 1.667499424E9, 1.667499472E9, 1.66749952E9, 1.667499568E9, 1.667499616E9, 1.667499664E9, 1.667499712E9, 1.66749976E9, 1.667499808E9, 1.667499856E9, 1.667499904E9, 1.667499952E9, 1.6675E9, 1.667500048E9, 1.667500096E9, 1.667500144E9, 1.667500192E9, 1.66750024E9, 1.66750056E9, 1.66750074E9, 1.667506564E9, 1.667506612E9, 1.66750666E9, 1.667506708E9, 1.667506756E9, 1.667506804E9, 1.667506852E9, 1.6675069E9, 1.667506948E9, 1.667506996E9, 1.667507044E9, 1.667507092E9, 1.66750714E9, 1.667507188E9, 1.667507236E9, 1.667507284E9, 1.667507332E9, 1.66750738E9, 1.667507428E9, 1.667507476E9, 1.667507524E9, 1.667507572E9, 1.66750762E9, 1.667507668E9, 1.667507716E9, 1.667507764E9, 1.667507812E9, 1.66750786E9, 1.667507908E9, 1.667507956E9, 1.667508004E9, 1.667508052E9, 1.6675081E9, 1.667508148E9, 1.667508196E9, 1.667508244E9, 1.667508292E9, 1.66750834E9, 1.667508388E9, 1.667508436E9, 1.667508484E9, 1.667508532E9, 1.66750858E9, 1.667508628E9, 1.667508676E9, 1.667508724E9, 1.667508772E9, 1.66750882E9, 1.667508868E9, 1.667508916E9, 1.667508964E9, 1.667509012E9, 1.66750906E9, 1.667509108E9, 1.667509156E9, 1.667509204E9, 1.667509252E9, 1.6675093E9, 1.667509348E9, 1.667509396E9, 1.667509444E9, 1.667509492E9, 1.66750954E9, 1.667509588E9, 1.667509636E9, 1.667509684E9, 1.667509732E9, 1.66750978E9, 1.66751016E9, 1.66751028E9, 1.667515867E9, 1.667515915E9, 1.667515963E9, 1.667516011E9, 1.667516059E9, 1.667516107E9, 1.667516155E9, 1.667516203E9, 1.667516251E9, 1.667516299E9, 1.667516347E9, 1.667516395E9, 1.667516443E9, 1.667516491E9, 1.667516539E9, 1.667516587E9, 1.667516635E9, 1.667516683E9, 1.667516731E9, 1.667516779E9, 1.667516827E9, 1.667516875E9, 1.667516923E9, 1.667516971E9, 1.667517019E9, 1.667517067E9, 1.667517115E9, 1.667517163E9, 1.667517211E9, 1.667517259E9, 1.667517307E9, 1.667517355E9, 1.667517403E9, 1.667517451E9, 1.667517499E9, 1.667517547E9, 1.667517595E9, 1.667517643E9, 1.667517691E9, 1.667517739E9, 1.667517787E9, 1.667517835E9, 1.667517883E9, 1.667517931E9, 1.667517979E9, 1.667518027E9, 1.667518075E9, 1.667518123E9, 1.667518171E9, 1.667518219E9, 1.667518267E9, 1.667518315E9, 1.667518363E9, 1.667518411E9, 1.667518459E9, 1.667518507E9, 1.667518555E9, 1.667518603E9, 1.667518651E9, 1.667518699E9, 1.667518747E9, 1.667518795E9, 1.667518843E9, 1.667518891E9, 1.667518939E9, 1.667518987E9, 1.667519035E9, 1.667519083E9, 1.667519131E9, 1.667519179E9, 1.66751952E9, 1.6675197E9, 1.667525152E9, 1.6675252E9, 1.667525248E9, 1.667525296E9, 1.667525344E9, 1.667525392E9, 1.66752544E9, 1.667525488E9, 1.667525536E9, 1.667525584E9, 1.667525632E9, 1.66752568E9, 1.667525728E9, 1.667525776E9, 1.667525824E9, 1.667525872E9, 1.66752592E9, 1.667525968E9, 1.667526016E9, 1.667526064E9, 1.667526112E9, 1.66752616E9, 1.667526208E9, 1.667526256E9, 1.667526304E9, 1.667526352E9, 1.6675264E9, 1.667526448E9, 1.667526496E9, 1.667526544E9, 1.667526592E9, 1.66752664E9, 1.667526688E9, 1.667526736E9, 1.667526784E9, 1.667526832E9, 1.66752688E9, 1.667526928E9, 1.667526976E9, 1.667527024E9, 1.667527072E9, 1.66752712E9, 1.667527168E9, 1.667527216E9, 1.667527264E9, 1.667527312E9, 1.66752736E9, 1.667527408E9, 1.667527456E9, 1.667527504E9, 1.667527552E9, 1.6675276E9, 1.667527648E9, 1.667527696E9, 1.667527744E9, 1.667527792E9, 1.66752784E9, 1.667527888E9, 1.667527936E9, 1.667527984E9, 1.667528032E9, 1.66752808E9, 1.667528128E9, 1.667528176E9, 1.667528224E9, 1.667528272E9, 1.66752832E9, 1.6675287E9, 1.66752894E9, 1.667534647E9, 1.667534695E9, 1.667534743E9, 1.667534791E9, 1.667534839E9, 1.667534887E9, 1.667534935E9, 1.667534983E9, 1.667535031E9, 1.667535079E9, 1.667535127E9, 1.667535175E9, 1.667535223E9, 1.667535271E9, 1.667535319E9, 1.667535367E9, 1.667535415E9, 1.667535463E9, 1.667535511E9, 1.667535559E9, 1.667535607E9, 1.667535655E9, 1.667535703E9, 1.667535751E9, 1.667535799E9, 1.667535847E9, 1.667535895E9, 1.667535943E9, 1.667535991E9, 1.667536039E9, 1.667536087E9, 1.667536135E9, 1.667536183E9, 1.667536231E9, 1.667536279E9, 1.667536327E9, 1.667536375E9, 1.667536423E9, 1.667536471E9, 1.667536519E9, 1.667536567E9, 1.667536615E9, 1.667536663E9, 1.667536711E9, 1.667536759E9, 1.667536807E9, 1.667536855E9, 1.667536903E9, 1.667536951E9, 1.667536999E9, 1.667537047E9, 1.667537095E9, 1.667537143E9, 1.667537191E9, 1.667537239E9, 1.667537287E9, 1.667537335E9, 1.667537383E9, 1.667537431E9, 1.667537479E9, 1.667537527E9, 1.667537575E9, 1.667537623E9, 1.667537671E9, 1.667537719E9, 1.667537767E9, 1.667537815E9, 1.667537863E9, 1.667537911E9, 1.667537959E9, 1.66753824E9, 1.66753842E9, 1.667544105E9, 1.667544153E9, 1.667544201E9, 1.667544249E9, 1.667544297E9, 1.667544345E9, 1.667544393E9, 1.667544441E9, 1.667544489E9, 1.667544537E9, 1.667544585E9, 1.667544633E9, 1.667544681E9, 1.667544729E9, 1.667544777E9, 1.667544825E9, 1.667544873E9, 1.667544921E9, 1.667544969E9, 1.667545017E9, 1.667545065E9, 1.667545113E9, 1.667545161E9, 1.667545209E9, 1.667545257E9, 1.667545305E9, 1.667545353E9, 1.667545401E9, 1.667545449E9, 1.667545497E9, 1.667545545E9, 1.667545593E9, 1.667545641E9, 1.667545689E9, 1.667545737E9, 1.667545785E9, 1.667545833E9, 1.667545881E9, 1.667545929E9, 1.667545977E9, 1.667546025E9, 1.667546073E9, 1.667546121E9, 1.667546169E9, 1.667546217E9, 1.667546265E9, 1.667546313E9, 1.667546361E9, 1.667546409E9, 1.667546457E9, 1.667546505E9, 1.667546553E9, 1.667546601E9, 1.667546649E9, 1.667546697E9, 1.667546745E9, 1.667546793E9, 1.667546841E9, 1.667546889E9, 1.667546937E9, 1.667546985E9, 1.667547033E9, 1.667547081E9, 1.667547129E9, 1.667547177E9, 1.667547225E9, 1.667547273E9, 1.667547321E9, 1.667547369E9, 1.66754772E9, 1.6675479E9, 1.667553492E9, 1.66755354E9, 1.667553588E9, 1.667553636E9, 1.667553684E9, 1.667553732E9, 1.66755378E9, 1.667553828E9, 1.667553876E9, 1.667553924E9, 1.667553972E9, 1.66755402E9, 1.667554068E9, 1.667554116E9, 1.667554164E9, 1.667554212E9, 1.66755426E9, 1.667554308E9, 1.667554356E9, 1.667554404E9, 1.667554452E9, 1.6675545E9, 1.667554548E9, 1.667554596E9, 1.667554644E9, 1.667554692E9, 1.66755474E9, 1.667554788E9, 1.667554836E9, 1.667554884E9, 1.667554932E9, 1.66755498E9, 1.667555028E9, 1.667555076E9, 1.667555124E9, 1.667555172E9, 1.66755522E9, 1.667555268E9, 1.667555316E9, 1.667555364E9, 1.667555412E9, 1.66755546E9, 1.667555508E9, 1.667555556E9, 1.667555604E9, 1.667555652E9, 1.6675557E9, 1.667555748E9, 1.667555796E9, 1.667555844E9, 1.667555892E9, 1.66755594E9, 1.667555988E9, 1.667556036E9, 1.667556084E9, 1.667556132E9, 1.66755618E9, 1.667556228E9, 1.667556276E9, 1.667556324E9, 1.667556372E9, 1.66755642E9, 1.667556468E9, 1.667556516E9, 1.667556564E9, 1.667556612E9, 1.66755666E9, 1.667556708E9, 1.667556756E9, 1.667556804E9, 1.667556852E9, 1.6675569E9, 1.66755726E9, 1.66755744E9, 1.667563171E9, 1.667563219E9, 1.667563267E9, 1.667563315E9, 1.667563363E9, 1.667563411E9, 1.667563459E9, 1.667563507E9, 1.667563555E9, 1.667563603E9, 1.667563651E9, 1.667563699E9, 1.667563747E9, 1.667563795E9, 1.667563843E9, 1.667563891E9, 1.667563939E9, 1.667563987E9, 1.667564035E9, 1.667564083E9, 1.667564131E9, 1.667564179E9, 1.667564227E9, 1.667564275E9, 1.667564323E9, 1.667564371E9, 1.667564419E9, 1.667564467E9, 1.667564515E9, 1.667564563E9, 1.667564611E9, 1.667564659E9, 1.667564707E9, 1.667564755E9, 1.667564803E9, 1.667564851E9, 1.667564899E9, 1.667564947E9, 1.667564995E9, 1.667565043E9, 1.667565091E9, 1.667565139E9, 1.667565187E9, 1.667565235E9, 1.667565283E9, 1.667565331E9, 1.667565379E9, 1.667565427E9, 1.667565475E9, 1.667565523E9, 1.667565571E9, 1.667565619E9, 1.667565667E9, 1.667565715E9, 1.667565763E9, 1.667565811E9, 1.667565859E9, 1.667565907E9, 1.667565955E9, 1.667566003E9, 1.667566051E9, 1.667566099E9, 1.667566147E9, 1.667566195E9, 1.667566243E9, 1.667566291E9, 1.667566339E9, 1.66756662E9, 1.6675668E9, 1.667572468E9, 1.667572516E9, 1.667572564E9, 1.667572612E9, 1.66757266E9, 1.667572708E9, 1.667572756E9, 1.667572804E9, 1.667572852E9, 1.6675729E9, 1.667572948E9, 1.667572996E9, 1.667573044E9, 1.667573092E9, 1.66757314E9, 1.667573188E9, 1.667573236E9, 1.667573284E9, 1.667573332E9, 1.66757338E9, 1.667573428E9, 1.667573476E9, 1.667573524E9, 1.667573572E9, 1.66757362E9, 1.667573668E9, 1.667573716E9, 1.667573764E9, 1.667573812E9, 1.66757386E9, 1.667573908E9, 1.667573956E9, 1.667574004E9, 1.667574052E9, 1.6675741E9, 1.667574148E9, 1.667574196E9, 1.667574244E9, 1.667574292E9, 1.66757434E9, 1.667574388E9, 1.667574436E9, 1.667574484E9, 1.667574532E9, 1.66757458E9, 1.667574628E9, 1.667574676E9, 1.667574724E9, 1.667574772E9, 1.66757482E9, 1.667574868E9, 1.667574916E9, 1.667574964E9, 1.667575012E9, 1.66757506E9, 1.667575108E9, 1.667575156E9, 1.667575204E9, 1.667575252E9, 1.6675753E9, 1.667575348E9, 1.667575396E9, 1.667575444E9, 1.667575492E9, 1.66757554E9, 1.667575588E9, 1.667575636E9, 1.667575684E9, 1.667575732E9, 1.66757578E9, 1.66757616E9, 1.66757634E9, 1.667581918E9, 1.667581966E9, 1.667582014E9, 1.667582062E9, 1.66758211E9, 1.667582158E9, 1.667582206E9, 1.667582254E9, 1.667582302E9, 1.66758235E9, 1.667582398E9, 1.667582446E9, 1.667582494E9, 1.667582542E9, 1.66758259E9, 1.667582638E9, 1.667582686E9, 1.667582734E9, 1.667582782E9, 1.66758283E9, 1.667582878E9, 1.667582926E9, 1.667582974E9, 1.667583022E9, 1.66758307E9, 1.667583118E9, 1.667583166E9, 1.667583214E9, 1.667583262E9, 1.66758331E9, 1.667583358E9, 1.667583406E9, 1.667583454E9, 1.667583502E9, 1.66758355E9, 1.667583598E9, 1.667583646E9, 1.667583694E9, 1.667583742E9, 1.66758379E9, 1.667583838E9, 1.667583886E9, 1.667583934E9, 1.667583982E9, 1.66758403E9, 1.667584078E9, 1.667584126E9, 1.667584174E9, 1.667584222E9, 1.66758427E9, 1.667584318E9, 1.667584366E9, 1.667584414E9, 1.667584462E9, 1.66758451E9, 1.667584558E9, 1.667584606E9, 1.667584654E9, 1.667584702E9, 1.66758475E9, 1.667584798E9, 1.667584846E9, 1.667584894E9, 1.667584942E9, 1.66758499E9, 1.667585038E9, 1.667585086E9, 1.667585134E9, 1.667585182E9, 1.66758523E9, 1.66758558E9, 1.66758576E9, 1.667591371E9, 1.667591419E9, 1.667591467E9, 1.667591515E9, 1.667591563E9, 1.667591611E9, 1.667591659E9, 1.667591707E9, 1.667591755E9, 1.667591803E9, 1.667591851E9, 1.667591899E9, 1.667591947E9, 1.667591995E9, 1.667592043E9, 1.667592091E9, 1.667592139E9, 1.667592187E9, 1.667592235E9, 1.667592283E9, 1.667592331E9, 1.667592379E9, 1.667592427E9, 1.667592475E9, 1.667592523E9, 1.667592571E9, 1.667592619E9, 1.667592667E9, 1.667592715E9, 1.667592763E9, 1.667592811E9, 1.667592859E9, 1.667592907E9, 1.667592955E9, 1.667593003E9, 1.667593051E9, 1.667593099E9, 1.667593147E9, 1.667593195E9, 1.667593243E9, 1.667593291E9, 1.667593339E9, 1.667593387E9, 1.667593435E9, 1.667593483E9, 1.667593531E9, 1.667593579E9, 1.667593627E9, 1.667593675E9, 1.667593723E9, 1.667593771E9, 1.667593819E9, 1.667593867E9, 1.667593915E9, 1.667593963E9, 1.667594011E9, 1.667594059E9, 1.667594107E9, 1.667594155E9, 1.667594203E9, 1.667594251E9, 1.667594299E9, 1.667594347E9, 1.667594395E9, 1.667594443E9, 1.667594491E9, 1.667594539E9, 1.66759482E9, 1.66759494E9, 1.66760064E9, 1.667600688E9, 1.667600736E9, 1.667600784E9, 1.667600832E9, 1.66760088E9, 1.667600928E9, 1.667600976E9, 1.667601024E9, 1.667601072E9, 1.66760112E9, 1.667601168E9, 1.667601216E9, 1.667601264E9, 1.667601312E9, 1.66760136E9, 1.667601408E9, 1.667601456E9, 1.667601504E9, 1.667601552E9, 1.6676016E9, 1.667601648E9, 1.667601696E9, 1.667601744E9, 1.667601792E9, 1.66760184E9, 1.667601888E9, 1.667601936E9, 1.667601984E9, 1.667602032E9, 1.66760208E9, 1.667602128E9, 1.667602176E9, 1.667602224E9, 1.667602272E9, 1.66760232E9, 1.667602368E9, 1.667602416E9, 1.667602464E9, 1.667602512E9, 1.66760256E9, 1.667602608E9, 1.667602656E9, 1.667602704E9, 1.667602752E9, 1.6676028E9, 1.667602848E9, 1.667602896E9, 1.667602944E9, 1.667602992E9, 1.66760304E9, 1.667603088E9, 1.667603136E9, 1.667603184E9, 1.667603232E9, 1.66760328E9, 1.667603328E9, 1.667603376E9, 1.667603424E9, 1.667603472E9, 1.66760352E9, 1.667603568E9, 1.667603616E9, 1.667603664E9, 1.667603712E9, 1.66760376E9, 1.667603808E9, 1.667603856E9, 1.667603904E9, 1.667603952E9, 1.667604E9, 1.6676043E9, 1.66760448E9, 1.667610334E9, 1.667610382E9, 1.66761043E9, 1.667610478E9, 1.667610526E9, 1.667610574E9, 1.667610622E9, 1.66761067E9, 1.667610718E9, 1.667610766E9, 1.667610814E9, 1.667610862E9, 1.66761091E9, 1.667610958E9, 1.667611006E9, 1.667611054E9, 1.667611102E9, 1.66761115E9, 1.667611198E9, 1.667611246E9, 1.667611294E9, 1.667611342E9, 1.66761139E9, 1.667611438E9, 1.667611486E9, 1.667611534E9, 1.667611582E9, 1.66761163E9, 1.667611678E9, 1.667611726E9, 1.667611774E9, 1.667611822E9, 1.66761187E9, 1.667611918E9, 1.667611966E9, 1.667612014E9, 1.667612062E9, 1.66761211E9, 1.667612158E9, 1.667612206E9, 1.667612254E9, 1.667612302E9, 1.66761235E9, 1.667612398E9, 1.667612446E9, 1.667612494E9, 1.667612542E9, 1.66761259E9, 1.667612638E9, 1.667612686E9, 1.667612734E9, 1.667612782E9, 1.66761283E9, 1.667612878E9, 1.667612926E9, 1.667612974E9, 1.667613022E9, 1.66761307E9, 1.667613118E9, 1.667613166E9, 1.667613214E9, 1.667613262E9, 1.66761331E9, 1.667613358E9, 1.667613406E9, 1.667613454E9, 1.667613502E9, 1.66761355E9, 1.667613598E9, 1.667613646E9, 1.667613694E9, 1.667613742E9, 1.66761379E9, 1.66761414E9, 1.66761432E9, 1.667620017E9, 1.667620065E9, 1.667620113E9, 1.667620161E9, 1.667620209E9, 1.667620257E9, 1.667620305E9, 1.667620353E9, 1.667620401E9, 1.667620449E9, 1.667620497E9, 1.667620545E9, 1.667620593E9, 1.667620641E9, 1.667620689E9, 1.667620737E9, 1.667620785E9, 1.667620833E9, 1.667620881E9, 1.667620929E9, 1.667620977E9, 1.667621025E9, 1.667621073E9, 1.667621121E9, 1.667621169E9, 1.667621217E9, 1.667621265E9, 1.667621313E9, 1.667621361E9, 1.667621409E9, 1.667621457E9, 1.667621505E9, 1.667621553E9, 1.667621601E9, 1.667621649E9, 1.667621697E9, 1.667621745E9, 1.667621793E9, 1.667621841E9, 1.667621889E9, 1.667621937E9, 1.667621985E9, 1.667622033E9, 1.667622081E9, 1.667622129E9, 1.667622177E9, 1.667622225E9, 1.667622273E9, 1.667622321E9, 1.667622369E9, 1.667622417E9, 1.667622465E9, 1.667622513E9, 1.667622561E9, 1.667622609E9, 1.667622657E9, 1.667622705E9, 1.667622753E9, 1.667622801E9, 1.667622849E9, 1.667622897E9, 1.667622945E9, 1.667622993E9, 1.667623041E9, 1.667623089E9, 1.667623137E9, 1.667623185E9, 1.667623233E9, 1.667623281E9, 1.667623329E9, 1.66762362E9, 1.6676238E9, 1.667629451E9, 1.667629499E9, 1.667629547E9, 1.667629595E9, 1.667629643E9, 1.667629691E9, 1.667629739E9, 1.667629787E9, 1.667629835E9, 1.667629883E9, 1.667629931E9, 1.667629979E9, 1.667630027E9, 1.667630075E9, 1.667630123E9, 1.667630171E9, 1.667630219E9, 1.667630267E9, 1.667630315E9, 1.667630363E9, 1.667630411E9, 1.667630459E9, 1.667630507E9, 1.667630555E9, 1.667630603E9, 1.667630651E9, 1.667630699E9, 1.667630747E9, 1.667630795E9, 1.667630843E9, 1.667630891E9, 1.667630939E9, 1.667630987E9, 1.667631035E9, 1.667631083E9, 1.667631131E9, 1.667631179E9, 1.667631227E9, 1.667631275E9, 1.667631323E9, 1.667631371E9, 1.667631419E9, 1.667631467E9, 1.667631515E9, 1.667631563E9, 1.667631611E9, 1.667631659E9, 1.667631707E9, 1.667631755E9, 1.667631803E9, 1.667631851E9, 1.667631899E9, 1.667631947E9, 1.667631995E9, 1.667632043E9, 1.667632091E9, 1.667632139E9, 1.667632187E9, 1.667632235E9, 1.667632283E9, 1.667632331E9, 1.667632379E9, 1.667632427E9, 1.667632475E9, 1.667632523E9, 1.667632571E9, 1.667632619E9, 1.66763292E9, 1.6676331E9, 1.667638814E9, 1.667638862E9, 1.66763891E9, 1.667638958E9, 1.667639006E9, 1.667639054E9, 1.667639102E9, 1.66763915E9, 1.667639198E9, 1.667639246E9, 1.667639294E9, 1.667639342E9, 1.66763939E9, 1.667639438E9, 1.667639486E9, 1.667639534E9, 1.667639582E9, 1.66763963E9, 1.667639678E9, 1.667639726E9, 1.667639774E9, 1.667639822E9, 1.66763987E9, 1.667639918E9, 1.667639966E9, 1.667640014E9, 1.667640062E9, 1.66764011E9, 1.667640158E9, 1.667640206E9, 1.667640254E9, 1.667640302E9, 1.66764035E9, 1.667640398E9, 1.667640446E9, 1.667640494E9, 1.667640542E9, 1.66764059E9, 1.667640638E9, 1.667640686E9, 1.667640734E9, 1.667640782E9, 1.66764083E9, 1.667640878E9, 1.667640926E9, 1.667640974E9, 1.667641022E9, 1.66764107E9, 1.667641118E9, 1.667641166E9, 1.667641214E9, 1.667641262E9, 1.66764131E9, 1.667641358E9, 1.667641406E9, 1.667641454E9, 1.667641502E9, 1.66764155E9, 1.667641598E9, 1.667641646E9, 1.667641694E9, 1.667641742E9, 1.66764179E9, 1.667641838E9, 1.667641886E9, 1.667641934E9, 1.667641982E9, 1.66764203E9, 1.66764234E9, 1.66764252E9, 1.667648246E9, 1.667648294E9, 1.667648342E9, 1.66764839E9, 1.667648438E9, 1.667648486E9, 1.667648534E9, 1.667648582E9, 1.66764863E9, 1.667648678E9, 1.667648726E9, 1.667648774E9, 1.667648822E9, 1.66764887E9, 1.667648918E9, 1.667648966E9, 1.667649014E9, 1.667649062E9, 1.66764911E9, 1.667649158E9, 1.667649206E9, 1.667649254E9, 1.667649302E9, 1.66764935E9, 1.667649398E9, 1.667649446E9, 1.667649494E9, 1.667649542E9, 1.66764959E9, 1.667649638E9, 1.667649686E9, 1.667649734E9, 1.667649782E9, 1.66764983E9, 1.667649878E9, 1.667649926E9, 1.667649974E9, 1.667650022E9, 1.66765007E9, 1.667650118E9, 1.667650166E9, 1.667650214E9, 1.667650262E9, 1.66765031E9, 1.667650358E9, 1.667650406E9, 1.667650454E9, 1.667650502E9, 1.66765055E9, 1.667650598E9, 1.667650646E9, 1.667650694E9, 1.667650742E9, 1.66765079E9, 1.667650838E9, 1.667650886E9, 1.667650934E9, 1.667650982E9, 1.66765103E9, 1.667651078E9, 1.667651126E9, 1.667651174E9, 1.667651222E9, 1.66765127E9, 1.667651318E9, 1.667651366E9, 1.667651414E9, 1.667651462E9, 1.66765151E9, 1.66765188E9, 1.667652E9, 1.667657672E9, 1.66765772E9, 1.667657768E9, 1.667657816E9, 1.667657864E9, 1.667657912E9, 1.66765796E9, 1.667658008E9, 1.667658056E9, 1.667658104E9, 1.667658152E9, 1.6676582E9, 1.667658248E9, 1.667658296E9, 1.667658344E9, 1.667658392E9, 1.66765844E9, 1.667658488E9, 1.667658536E9, 1.667658584E9, 1.667658632E9, 1.66765868E9, 1.667658728E9, 1.667658776E9, 1.667658824E9, 1.667658872E9, 1.66765892E9, 1.667658968E9, 1.667659016E9, 1.667659064E9, 1.667659112E9, 1.66765916E9, 1.667659208E9, 1.667659256E9, 1.667659304E9, 1.667659352E9, 1.6676594E9, 1.667659448E9, 1.667659496E9, 1.667659544E9, 1.667659592E9, 1.66765964E9, 1.667659688E9, 1.667659736E9, 1.667659784E9, 1.667659832E9, 1.66765988E9, 1.667659928E9, 1.667659976E9, 1.667660024E9, 1.667660072E9, 1.66766012E9, 1.667660168E9, 1.667660216E9, 1.667660264E9, 1.667660312E9, 1.66766036E9, 1.667660408E9, 1.667660456E9, 1.667660504E9, 1.667660552E9, 1.6676606E9, 1.667660648E9, 1.667660696E9, 1.667660744E9, 1.667660792E9, 1.66766084E9, 1.667660888E9, 1.667660936E9, 1.667660984E9, 1.667661032E9, 1.66766108E9, 1.66766136E9, 1.66766154E9, 1.667667297E9, 1.667667345E9, 1.667667393E9, 1.667667441E9, 1.667667489E9, 1.667667537E9, 1.667667585E9, 1.667667633E9, 1.667667681E9, 1.667667729E9, 1.667667777E9, 1.667667825E9, 1.667667873E9, 1.667667921E9, 1.667667969E9, 1.667668017E9, 1.667668065E9, 1.667668113E9, 1.667668161E9, 1.667668209E9, 1.667668257E9, 1.667668305E9, 1.667668353E9, 1.667668401E9, 1.667668449E9, 1.667668497E9, 1.667668545E9, 1.667668593E9, 1.667668641E9, 1.667668689E9, 1.667668737E9, 1.667668785E9, 1.667668833E9, 1.667668881E9, 1.667668929E9, 1.667668977E9, 1.667669025E9, 1.667669073E9, 1.667669121E9, 1.667669169E9, 1.667669217E9, 1.667669265E9, 1.667669313E9, 1.667669361E9, 1.667669409E9, 1.667669457E9, 1.667669505E9, 1.667669553E9, 1.667669601E9, 1.667669649E9, 1.667669697E9, 1.667669745E9, 1.667669793E9, 1.667669841E9, 1.667669889E9, 1.667669937E9, 1.667669985E9, 1.667670033E9, 1.667670081E9, 1.667670129E9, 1.667670177E9, 1.667670225E9, 1.667670273E9, 1.667670321E9, 1.667670369E9, 1.667670417E9, 1.667670465E9, 1.667670513E9, 1.667670561E9, 1.667670609E9, 1.6676709E9, 1.66767108E9, 1.667676687E9, 1.667676735E9, 1.667676783E9, 1.667676831E9, 1.667676879E9, 1.667676927E9, 1.667676975E9, 1.667677023E9, 1.667677071E9, 1.667677119E9, 1.667677167E9, 1.667677215E9, 1.667677263E9, 1.667677311E9, 1.667677359E9, 1.667677407E9, 1.667677455E9, 1.667677503E9, 1.667677551E9, 1.667677599E9, 1.667677647E9, 1.667677695E9, 1.667677743E9, 1.667677791E9, 1.667677839E9, 1.667677887E9, 1.667677935E9, 1.667677983E9, 1.667678031E9, 1.667678079E9, 1.667678127E9, 1.667678175E9, 1.667678223E9, 1.667678271E9, 1.667678319E9, 1.667678367E9, 1.667678415E9, 1.667678463E9, 1.667678511E9, 1.667678559E9, 1.667678607E9, 1.667678655E9, 1.667678703E9, 1.667678751E9, 1.667678799E9, 1.667678847E9, 1.667678895E9, 1.667678943E9, 1.667678991E9, 1.667679039E9, 1.667679087E9, 1.667679135E9, 1.667679183E9, 1.667679231E9, 1.667679279E9, 1.667679327E9, 1.667679375E9, 1.667679423E9, 1.667679471E9, 1.667679519E9, 1.667679567E9, 1.667679615E9, 1.667679663E9, 1.667679711E9, 1.667679759E9, 1.667679807E9, 1.667679855E9, 1.667679903E9, 1.667679951E9, 1.667679999E9, 1.66768038E9, 1.66768056E9, 1.667686333E9, 1.667686381E9, 1.667686429E9, 1.667686477E9, 1.667686525E9, 1.667686573E9, 1.667686621E9, 1.667686669E9, 1.667686717E9, 1.667686765E9, 1.667686813E9, 1.667686861E9, 1.667686909E9, 1.667686957E9, 1.667687005E9, 1.667687053E9, 1.667687101E9, 1.667687149E9, 1.667687197E9, 1.667687245E9, 1.667687293E9, 1.667687341E9, 1.667687389E9, 1.667687437E9, 1.667687485E9, 1.667687533E9, 1.667687581E9, 1.667687629E9, 1.667687677E9, 1.667687725E9, 1.667687773E9, 1.667687821E9, 1.667687869E9, 1.667687917E9, 1.667687965E9, 1.667688013E9, 1.667688061E9, 1.667688109E9, 1.667688157E9, 1.667688205E9, 1.667688253E9, 1.667688301E9, 1.667688349E9, 1.667688397E9, 1.667688445E9, 1.667688493E9, 1.667688541E9, 1.667688589E9, 1.667688637E9, 1.667688685E9, 1.667688733E9, 1.667688781E9, 1.667688829E9, 1.667688877E9, 1.667688925E9, 1.667688973E9, 1.667689021E9, 1.667689069E9, 1.667689117E9, 1.667689165E9, 1.667689213E9, 1.667689261E9, 1.667689309E9, 1.667689357E9, 1.667689405E9, 1.667689453E9, 1.667689501E9, 1.667689549E9, 1.6676898E9}
    LATITUDE = 
      {37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4165, 37.4383, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4385, 37.4525, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4527, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4642, 37.4762, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.476, 37.4847, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.4843, 37.488, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.4878, 37.49, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4897, 37.4948, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4945, 37.4987, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.4982, 37.5023, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.5015, 37.4985, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.4978, 37.493, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4918, 37.4888, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.488, 37.4918, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4912, 37.4958, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.4957, 37.496, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4962, 37.4992, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.499, 37.5035, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.5032, 37.509, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5087, 37.5093, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.5092, 37.508, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5073, 37.5087, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5083, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.5175, 37.524, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5237, 37.5267, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.526, 37.5288, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5282, 37.5348, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5343, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5423, 37.5515, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.552, 37.5593, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5598, 37.5635, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5638, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.5722, 37.584, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5838, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.5942, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6037, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6135, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6267, 37.6417, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6418, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.6522, 37.661, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.6608, 37.673, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6727, 37.6923, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.692, 37.7083, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7082, 37.7202, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7203, 37.7317, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7318, 37.7455, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7453, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7605, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7747, 37.7852, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.785, 37.798, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.7978, 37.8133, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8135, 37.8273, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8275, 37.8373, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.837, 37.8443, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.844, 37.857, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8563, 37.8728, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8727, 37.8862, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.886, 37.8948, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.8945, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9033, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9178, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9368, 37.9503, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9505, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9585, 37.9695}
    LONGITUDE = 
      {-126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -126.0032, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9858, -125.9623, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9625, -125.9347, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9348, -125.9088, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.9092, -125.8858, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8867, -125.8582, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8592, -125.8303, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8308, -125.8092, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.8098, -125.7898, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.7908, -125.774, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7748, -125.7555, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7558, -125.7413, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7415, -125.7318, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7327, -125.7292, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7305, -125.7232, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7238, -125.7083, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.7088, -125.6978, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6982, -125.6907, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.691, -125.6828, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.6832, -125.67, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6705, -125.6578, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6582, -125.6512, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6518, -125.6473, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6477, -125.6337, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6342, -125.6187, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6192, -125.6025, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.6032, -125.5942, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.595, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.5853, -125.569, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5695, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5475, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.5183, -125.4938, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4935, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4712, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.4495, -125.425, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.4253, -125.3993, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3992, -125.3705, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3707, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3395, -125.3012, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.301, -125.2605, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.26, -125.2253, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.225, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1948, -125.1592, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1595, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.1188, -125.0763, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0758, -125.0393, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0388, -125.0087, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -125.0082, -124.976, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9758, -124.9457, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.9455, -124.915, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.9152, -124.8817, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.8815, -124.846, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8457, -124.8135, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.8133, -124.7847, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7843, -124.7602, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7598, -124.7333, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7335, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.7037, -124.6717, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.6712, -124.64, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.6397, -124.609, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.6085, -124.5815, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5812, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5492, -124.5177, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.5173, -124.4875}
    DEPTH = 
      {NaN, 500.27908, 495.76392, 489.58514, 481.34647, 473.34512, 465.50192, 457.3415, 449.18076, 441.17816, 433.413, 425.64752, 417.88174, 410.35342, 402.98334, 395.29596, 387.6083, 379.8411, 371.75656, 363.59244, 355.26944, 347.10468, 338.62247, 330.45703, 322.2913, 314.20447, 306.27594, 298.2678, 290.10074, 282.0127, 273.845, 265.7563, 257.66727, 249.65724, 241.6469, 233.55693, 225.70459, 217.77263, 210.07834, 202.38377, 195.00623, 187.66808, 180.29, 173.229, 166.24712, 159.34433, 152.28262, 145.14133, 137.76172, 130.61992, 123.55722, 116.653, 110.542175, 104.3518, 98.08187, 92.129234, 86.097046, 80.38219, 74.74654, 68.8726, 62.601585, 56.092228, 49.74144, 43.54923, 37.912567, 32.593323, 27.750305, 23.224762, 18.699118, 14.093973, 8.615305, 3.4541059, NaN, NaN, 501.2289, 496.71378, 490.69345, 482.21716, 473.2652, 463.8375, 454.33014, 444.82233, 435.23483, 425.4884, 415.97928, 406.4697, 397.19745, 387.84552, 378.81018, 369.93298, 361.05542, 352.65308, 344.2504, 335.60953, 327.20615, 318.961, 310.95337, 302.78683, 294.69928, 286.5321, 278.52322, 270.6726, 262.6631, 254.49466, 246.4052, 238.31543, 230.62192, 222.8488, 215.15471, 207.46034, 199.76567, 192.46738, 185.16881, 177.79065, 170.61058, 163.54927, 156.56706, 149.34657, 142.36388, 135.1429, 128.08037, 121.17631, 113.795845, 105.85957, 98.31983, 90.70044, 83.23952, 76.96895, 71.65073, 66.09423, 60.22005, 54.10755, 48.074253, 42.19956, 36.602562, 31.600864, 26.916622, 21.517702, 15.801042, 9.607814, 3.414399, NaN, NaN, 501.5848, 497.30734, 491.5247, 483.6822, 476.15628, 468.31323, 460.46985, 452.3885, 444.3068, 436.22482, 427.82553, 419.7429, 411.50146, 403.49744, 395.41382, 387.0129, 378.4531, 369.97223, 361.491, 353.2472, 344.8842, 336.4812, 328.3157, 320.0706, 311.5873, 303.5001, 295.41257, 287.40405, 279.39517, 270.59302, 262.1077, 253.93922, 246.167, 238.31517, 230.62167, 222.68993, 215.07515, 207.46011, 200.00343, 192.5465, 185.6446, 178.58382, 172.07817, 165.25493, 158.51082, 151.6078, 144.30779, 137.48364, 130.57991, 123.43787, 116.4543, 109.073685, 102.08963, 95.58154, 88.75577, 82.08852, 75.34167, 68.75336, 62.323593, 56.290546, 50.3764, 44.343, 39.023933, 33.466557, 28.067814, 22.510136, 16.475916, 11.314928, 6.2332134, 2.34244, NaN, NaN, 501.78232, 497.3464, 491.3261, 483.00833, 474.7694, 466.45093, 457.57755, 448.8622, 440.305, 431.58896, 422.3971, 413.44254, 404.09137, 394.8983, 385.86328, 376.66937, 367.31653, 358.28033, 349.16446, 340.9202, 332.63596, 324.1532, 315.90793, 307.9002, 299.57498, 290.93228, 282.5271, 273.40787, 264.05032, 255.08891, 245.96848, 237.48213, 228.75749, 220.5084, 212.02101, 203.85059, 195.67982, 187.11208, 178.70264, 170.76889, 163.0332, 155.09885, 147.16418, 139.38792, 131.92879, 124.23131, 116.37482, 108.9942, 101.53396, 94.54965, 87.644485, 81.05657, 74.46845, 67.48322, 60.577137, 54.06774, 47.875683, 41.842216, 35.411617, 29.29839, 24.137732, 18.579954, 13.419024, 8.257965, 4.0496206, NaN, NaN, 500.07886, 495.6429, 489.781, 481.2255, 472.82806, 463.95496, 455.2399, 446.84143, 438.6803, 430.51886, 422.43634, 414.512, 406.27036, 398.26614, 390.18237, 382.09827, 374.0931, 366.4047, 358.55746, 350.70993, 342.78284, 334.69687, 326.6106, 318.60327, 310.43707, 301.8741, 293.3901, 284.82642, 276.1038, 267.2222, 258.49884, 249.6958, 240.73375, 232.00925, 222.8878, 214.40051, 205.91287, 197.58356, 189.65054, 181.8759, 174.10095, 166.64308, 159.1056, 151.72653, 144.50589, 137.52306, 130.38127, 123.39796, 116.57312, 109.66869, 103.160866, 96.652824, 89.27151, 82.52491, 75.77809, 69.50732, 63.553875, 57.44149, 51.725853, 45.53373, 38.745995, 32.87105, 27.392908, 22.390999, 17.230171, 12.069212, 6.431708, 2.4615417, NaN, NaN, 500.19745, 495.6823, 489.7412, 481.50256, 473.81815, 465.81656, 458.05234, 449.81244, 442.0476, 434.0448, 426.1209, 418.3552, 410.74768, 402.82288, 395.29404, 387.68567, 380.07703, 372.78516, 365.25522, 357.725, 350.2738, 342.42596, 334.6571, 326.88794, 319.19775, 311.34872, 303.658, 295.4119, 287.0069, 278.91876, 270.8303, 262.6622, 254.41449, 246.40437, 238.63187, 230.77977, 223.00668, 215.2333, 207.77693, 200.47894, 193.41869, 186.35818, 179.6941, 173.10916, 166.60335, 160.01799, 153.35306, 146.92596, 140.41931, 133.75375, 127.2467, 120.739426, 114.07323, 107.248085, 100.184616, 93.75585, 87.32689, 80.89773, 74.07148, 67.245, 60.81521, 54.623363, 48.510715, 42.39789, 36.60244, 31.600758, 26.837135, 22.311594, 17.468359, 12.307407, 6.90812, 2.6997528, NaN, NaN, 500.63303, 496.2763, 490.57288, 482.41348, 474.41223, 465.6184, 457.0619, 448.58426, 439.9478, 431.62796, 423.387, 415.06647, 406.7456, 398.4244, 390.02362, 381.86026, 373.69656, 365.61185, 357.6853, 349.59995, 341.4746, 333.0715, 324.8266, 316.42282, 308.57367, 300.64496, 292.71594, 284.7073, 276.53976, 268.60983, 261.07608, 253.70067, 246.48363, 239.66289, 232.60397, 225.62413, 218.4061, 211.26714, 203.7313, 196.67114, 189.49176, 182.27246, 174.89423, 167.27771, 159.6609, 152.04382, 144.10905, 136.25334, 128.63539, 120.93779, 113.319275, 105.70047, 97.922646, 90.70012, 83.715454, 77.04805, 70.301056, 64.03011, 57.52084, 51.170124, 44.819214, 38.547497, 32.59316, 27.035616, 21.716116, 16.634672, 11.553102, 6.3920026, 2.8188581, NaN, NaN, 501.38535, 496.71182, 490.6915, 483.08667, 475.56076, 467.48, 459.31973, 451.23834, 443.07742, 434.8369, 426.91306, 418.90964, 411.06442, 403.13965, 395.21457, 387.28918, 378.88794, 370.96194, 362.79782, 354.47485, 346.50827, 338.0261, 329.54355, 321.13995, 313.05316, 305.04532, 297.19577, 289.10803, 281.33716, 273.64526, 265.8738, 258.02277, 250.72656, 243.35078, 235.7368, 228.51913, 221.38052, 214.47963, 207.5785, 200.35983, 193.06158, 185.8424, 178.2263, 170.68924, 163.15192, 155.69365, 148.07643, 140.53827, 133.47595, 126.492744, 119.5093, 112.208176, 104.98615, 98.16071, 91.33504, 84.58852, 77.92114, 71.01543, 63.871334, 56.806374, 49.62209, 42.874195, 36.7612, 30.489237, 23.026146, 16.118574, 10.560589, 5.161258, 1.9851147, NaN, NaN, 498.65234, 493.97876, 487.72073, 478.76904, 470.21307, 461.736, 453.57547, 445.49387, 437.80814, 430.1221, 422.35654, 414.66995, 407.0623, 399.53363, 391.9254, 384.31696, 376.7082, 368.78207, 361.01422, 353.4046, 345.7947, 337.9467, 329.93982, 321.77408, 313.68732, 305.7588, 297.5921, 289.42508, 281.01987, 273.01077, 264.7635, 256.67447, 248.74376, 240.73343, 232.40552, 224.31523, 216.06598, 207.89572, 199.96312, 192.18887, 184.29533, 176.28249, 168.66603, 161.52534, 154.78113, 148.43344, 142.56165, 136.68968, 131.21432, 125.81817, 120.10445, 114.39056, 108.67651, 103.04168, 97.96226, 93.04144, 88.27926, 83.59633, 78.43705, 72.72201, 66.29239, 59.783188, 53.27378, 46.843555, 39.77801, 33.585533, 28.186813, 23.105534, 17.706535, 11.989795, 6.193492, 2.3821344, NaN, NaN, 500.43445, 495.84012, 489.74057, 481.10587, 472.70844, 463.7561, 455.04108, 446.32565, 437.76837, 429.6069, 421.28665, 413.20377, 405.04135, 396.87857, 388.87402, 381.02765, 373.1017, 365.09622, 356.6941, 348.29163, 339.65097, 331.08923, 322.05148, 313.25116, 304.2919, 295.17365, 285.89642, 276.5395, 267.1821, 257.6657, 248.4661, 239.26607, 229.907, 220.70615, 211.66353, 203.01715, 194.52905, 186.11995, 177.7105, 169.61806, 161.803, 154.42403, 147.20349, 140.22076, 133.15845, 126.17523, 119.19178, 112.04937, 104.82735, 98.081276, 91.73183, 85.144066, 78.238594, 71.571014, 65.141365, 58.711514, 52.678383, 46.96262, 40.84975, 34.57792, 28.583775, 23.264318, 17.944725, 12.148592, 6.2728925, 2.7791533, NaN, NaN, 499.56323, 494.96887, 488.94852, 480.9475, 473.02542, 464.78613, 456.62573, 448.46503, 440.1455, 431.98413, 423.82245, 415.81894, 407.8151, 399.49396, 390.9347, 382.61285, 374.21143, 365.80966, 357.40756, 348.68802, 340.16632, 331.52533, 323.04254, 314.16296, 305.5209, 296.79916, 288.15634, 279.59247, 271.02826, 262.38437, 254.13664, 245.49203, 237.085, 228.59833, 220.50789, 212.6551, 204.88135, 197.42459, 189.80893, 182.35164, 175.01308, 167.6346, 160.25584, 153.0355, 145.73558, 138.27669, 130.81754, 123.9136, 117.168144, 110.5812, 104.07341, 97.56541, 91.37468, 84.94565, 78.59579, 72.08698, 65.33983, 58.671833, 52.083008, 46.04968, 40.33373, 34.697014, 29.139534, 24.058279, 18.500513, 12.466194, 6.193491, 2.461538, NaN, NaN, 502.29623, 497.86038, 491.9193, 483.6808, 475.4419, 467.12347, 458.4878, 450.01022, 441.13614, 432.7371, 424.25845, 415.77948, 407.61716, 399.53375, 391.37076, 383.1282, 374.96457, 366.6421, 358.24002, 349.8376, 341.55374, 333.15063, 324.7472, 316.3434, 307.62213, 299.13834, 290.6542, 282.32834, 274.0814, 266.07205, 258.30032, 250.21104, 242.28008, 234.74536, 227.2897, 219.75446, 212.4569, 205.07974, 197.623, 190.32466, 182.94672, 175.88586, 168.82477, 161.76341, 154.46379, 147.32262, 140.10182, 132.72208, 125.34207, 117.72372, 110.501884, 103.67663, 97.08925, 90.581024, 84.15196, 78.119576, 72.08701, 66.21303, 60.2595, 53.988255, 47.875595, 41.603973, 35.570335, 29.774696, 23.8995, 18.659317, 13.2602, 7.860941, 3.652596, NaN, NaN, 501.62317, 497.26648, 491.40463, 483.64136, 476.27393, 468.58932, 460.74597, 453.0608, 445.61304, 437.61035, 429.2904, 421.44556, 413.6797, 405.83426, 397.90927, 389.82547, 381.89987, 373.65695, 365.25516, 357.01154, 348.80722, 340.64224, 332.47693, 324.46985, 316.62103, 308.8512, 301.08105, 293.38992, 286.09497, 278.64117, 271.2664, 263.97064, 256.75397, 249.45772, 242.24051, 234.86444, 227.4881, 220.27013, 213.13123, 205.83342, 198.6147, 191.3957, 184.17647, 177.03632, 169.81657, 162.59657, 155.45567, 148.15582, 140.69702, 133.23793, 125.937294, 118.16024, 109.98608, 101.73222, 93.47804, 85.302895, 77.76242, 70.38043, 63.474453, 57.04454, 50.93197, 45.057377, 39.658955, 34.260387, 28.385319, 22.589476, 16.15828, 9.488677, 3.9305098, NaN, NaN, 500.51413, 495.9198, 489.82025, 480.94788, 471.59976, 462.33047, 453.06076, 444.10754, 435.15396, 425.88303, 416.69092, 407.57767, 398.62247, 389.66693, 380.79022, 372.0717, 363.35275, 354.47495, 345.676, 337.03525, 328.55267, 320.46616, 312.30005, 304.37146, 296.44257, 288.4341, 280.5046, 272.9713, 265.7549, 258.6176, 251.71796, 244.8974, 238.15591, 231.65216, 225.14821, 218.80267, 212.45695, 206.11104, 199.60626, 193.18062, 186.67545, 180.17006, 173.26778, 166.36526, 159.30385, 152.16283, 144.78351, 137.24522, 129.4686, 121.69168, 113.59702, 105.422676, 97.486115, 89.94609, 82.326416, 75.18272, 68.197525, 61.370857, 54.067657, 47.002357, 40.730705, 35.17339, 29.61592, 24.37588, 19.69149, 14.1336, 7.622737, 3.0967712, NaN, NaN, 497.9792, 493.22635, 487.28516, 479.99707, 473.10483, 465.57858, 457.8936, 450.44598, 443.07736, 435.62924, 428.4978, 421.2869, 414.15497, 406.94354, 399.57336, 392.2029, 384.99072, 377.7783, 370.88263, 363.82822, 356.37723, 349.00525, 341.633, 334.33975, 326.96698, 319.59396, 312.69635, 305.71924, 298.74188, 291.28854, 283.99353, 276.53964, 269.0855, 261.63107, 254.2557, 246.56282, 238.86964, 231.49345, 224.03767, 216.58162, 209.40294, 202.26366, 194.88615, 187.66704, 180.36833, 173.06938, 165.77016, 158.39134, 150.85356, 143.63289, 136.65004, 129.50824, 122.207466, 114.74771, 107.12897, 99.66866, 92.049355, 84.42976, 77.36552, 69.74538, 62.918762, 56.09192, 49.97932, 44.34287, 39.1826, 33.942806, 28.147123, 21.080933, 14.729091, 8.456454, 3.0570683, NaN, NaN, 498.09793, 493.50354, 487.56238, 479.87817, 472.27295, 464.2713, 456.19012, 448.26706, 440.34372, 432.49933, 424.81308, 417.2058, 409.59827, 402.30743, 394.9371, 387.5665, 379.72006, 372.1904, 364.73972, 357.52658, 350.35278, 342.9806, 335.7667, 328.6318, 321.4174, 314.1234, 306.67065, 299.29688, 291.76425, 284.31067, 277.0154, 269.56128, 262.26547, 254.6522, 246.95934, 239.4248, 231.73137, 224.11697, 216.74023, 209.36325, 201.90666, 194.6878, 187.38936, 180.40799, 173.34705, 165.96849, 158.82771, 151.84537, 144.8628, 137.95932, 131.29369, 124.548485, 117.96178, 111.374855, 104.70835, 98.27974, 91.85092, 85.81876, 79.945175, 74.38892, 68.911896, 63.117207, 57.242966, 51.6861, 46.049694, 40.33374, 34.9352, 29.53651, 24.137682, 18.659313, 13.895395, 9.448972, 4.6054354, 1.9057101, NaN, NaN, 499.08798, 494.4144, 488.39404, 479.52158, 470.49033, 461.37943, 452.4266, 444.028, 435.3914, 426.83362, 418.19626, 409.55856, 401.2375, 392.83682, 384.35654, 376.19296, 367.712, 359.15146, 350.5905, 341.94998, 333.46762, 325.30203, 316.97754, 308.6527, 300.40686, 292.31924, 284.5485, 276.53955, 268.6889, 260.75867, 252.51086, 244.57999, 236.49019, 228.16211, 219.67505, 211.50494, 203.09653, 195.08441, 186.99265, 179.13858, 171.60156, 163.7469, 155.97128, 148.43343, 140.97462, 133.67427, 126.45301, 119.46957, 112.485886, 105.26388, 98.27972, 91.454056, 84.62817, 77.80205, 71.37259, 65.181076, 59.465656, 53.6707, 47.954964, 42.318455, 36.761185, 31.283154, 25.804977, 20.406052, 15.4833765, 10.084179, 4.8436437, 1.8263054, NaN, NaN, 501.0285, 496.75104, 491.1268, 482.65057, 473.85712, 465.14252, 456.586, 448.4253, 440.34348, 432.3406, 424.41666, 416.25464, 408.33008, 400.48447, 392.4008, 384.23752, 376.1532, 368.06857, 359.90436, 351.8191, 343.2975, 334.8152, 326.0947, 317.69098, 309.44547, 301.12036, 292.557, 284.3898, 275.82578, 267.57858, 259.4897, 251.24185, 242.83507, 234.34863, 226.09978, 217.92993, 209.36313, 201.03395, 192.70445, 184.1366, 175.72707, 167.31718, 158.9863, 150.81378, 142.56158, 134.30905, 126.373604, 118.675934, 111.37479, 104.15274, 97.00981, 89.946, 82.96132, 76.77015, 70.8963, 65.339806, 59.94193, 54.46452, 48.35188, 42.31844, 36.205437, 30.17164, 24.137669, 18.341711, 12.783791, 7.146317, 2.7791529, NaN, NaN, 501.1471, 496.55276, 490.53247, 481.81857, 472.7874, 463.9143, 455.04083, 446.2462, 437.60965, 428.97275, 421.52414, 413.20355, 404.88263, 396.3236, 387.68497, 378.96674, 370.7237, 362.79736, 354.87076, 346.94382, 338.85803, 331.08905, 323.31976, 315.6295, 307.85962, 300.08945, 292.5569, 285.10333, 277.5702, 270.0368, 262.82034, 255.5243, 248.06941, 241.09012, 234.11058, 227.05148, 220.2301, 213.09122, 205.95209, 198.73337, 191.3954, 183.93817, 176.56001, 169.1816, 161.88223, 154.58263, 146.64798, 139.03043, 131.25388, 123.39768, 115.46182, 107.68439, 100.065384, 92.4461, 85.4615, 78.39729, 71.88849, 65.61761, 59.584682, 53.630962, 47.67707, 41.802395, 36.086334, 30.449503, 24.733124, 19.334173, 14.411477, 8.932853, 3.7716968, NaN, NaN, 499.84003, 495.4041, 489.5422, 482.175, 474.96594, 467.36053, 459.6756, 451.91116, 444.3049, 436.3022, 428.53687, 420.6128, 413.00537, 405.55618, 397.9482, 390.49844, 383.1277, 375.75668, 368.3854, 361.01385, 353.44388, 346.15106, 338.38235, 330.69263, 323.08188, 315.55014, 307.78027, 300.01013, 292.2397, 284.46893, 276.7772, 269.00586, 261.63074, 254.33469, 247.19698, 239.82109, 232.8415, 225.8617, 219.04028, 212.13931, 205.43643, 198.53502, 191.4747, 184.89015, 178.22604, 171.48239, 164.57983, 157.5977, 150.29794, 142.75987, 134.90411, 127.286125, 119.74721, 111.96993, 104.35109, 97.28754, 90.38248, 83.7153, 77.52416, 71.57097, 65.81605, 60.180035, 54.464485, 48.828163, 43.191685, 36.99932, 30.965553, 25.328583, 19.770855, 14.609973, 9.607762, 4.129011, NaN, NaN, 501.3451, 496.83, 490.73047, 482.5711, 474.49066, 465.8553, 457.37805, 449.21735, 441.05637, 432.97427, 424.81262, 416.49216, 408.09213, 399.69174, 390.89474, 382.33514, 373.7752, 365.29416, 356.81277, 348.33102, 340.00748, 331.52505, 323.12155, 314.7177, 306.3135, 297.98828, 289.50412, 281.25748, 273.0898, 264.92184, 256.51562, 248.34697, 240.0987, 231.92941, 223.60115, 215.35188, 207.02295, 198.93167, 190.60208, 182.66882, 175.21127, 167.75346, 160.37473, 153.07506, 145.5371, 138.31625, 130.77774, 122.6041, 114.66821, 106.57329, 98.47805, 90.382484, 83.08033, 76.1748, 69.74529, 63.394966, 56.965065, 50.69373, 44.898525, 39.42072, 34.101547, 29.099815, 23.780376, 18.222605, 12.347084, 6.3125896, 2.1042182, NaN, NaN, 500.43414, 495.91904, 490.374, 482.37305, 474.45105, 466.4495, 458.28915, 450.1285, 442.20526, 434.1232, 425.9616, 417.72043, 409.3997, 401.15787, 392.5987, 383.88068, 375.71707, 367.2361, 358.91333, 350.74875, 342.3064, 333.9826, 325.65848, 317.25476, 309.3264, 301.08054, 292.91367, 284.5086, 276.02386, 267.6181, 259.2913, 251.04346, 243.11253, 235.2606, 227.24976, 219.31792, 211.22713, 203.37398, 195.3619, 187.34949, 179.41609, 171.40306, 163.46907, 155.53476, 147.67949, 140.06198, 132.52353, 125.22288, 118.08068, 110.93824, 103.79555, 97.12881, 90.69997, 84.27092, 77.92104, 71.17409, 64.42691, 57.44136, 50.931885, 44.977913, 39.10316, 33.307632, 27.511936, 22.11306, 16.237652, 10.520874, 5.2009525, 1.7071975, NaN, NaN, 501.42398, 497.06732, 491.28467, 483.0461, 474.88647, 466.25113, 457.53622, 448.7417, 440.26373, 432.1816, 423.86148, 415.46173, 407.1409, 398.26498, 389.38867, 380.43274, 371.55566, 362.75748, 354.03818, 345.08072, 336.4003, 327.91772, 319.5141, 311.03082, 302.86435, 294.93542, 287.08548, 279.15594, 271.46402, 263.8511, 256.3965, 248.78302, 241.08995, 233.39659, 225.70294, 217.53308, 209.28357, 201.03372, 192.3869, 183.97772, 176.00453, 168.30875, 160.77133, 153.313, 145.8544, 138.55423, 131.33315, 124.27052, 116.96958, 109.58901, 102.44628, 95.22393, 88.080696, 80.93721, 73.55534, 66.570114, 59.425877, 52.678318, 46.48624, 40.532146, 34.974834, 29.258583, 24.018547, 18.460787, 13.061676, 8.05943, 3.2952735, NaN, NaN, 499.79984, 495.2847, 489.26437, 480.94653, 472.78677, 464.5475, 455.99097, 447.59253, 439.1938, 430.79468, 422.39523, 414.2332, 405.99155, 397.9081, 389.7451, 381.2647, 372.784, 364.46143, 356.2971, 347.81534, 339.4918, 331.24716, 323.1608, 314.75696, 306.35278, 298.10684, 289.78128, 281.93115, 274.16, 265.9921, 258.45828, 251.0035, 243.38982, 236.17242, 228.71683, 220.62642, 212.69432, 204.3653, 196.1946, 188.26157, 180.44724, 172.67226, 165.05568, 157.51817, 150.5358, 143.3945, 136.09424, 129.26985, 122.60395, 116.01719, 109.27149, 102.76367, 96.335014, 89.82678, 83.79458, 77.60345, 71.41213, 65.37938, 58.94955, 52.83705, 47.041916, 41.484787, 35.9275, 30.37007, 24.73309, 19.413546, 14.0144615, 8.85344, 4.803932, 1.9454075, NaN, NaN, 499.87888, 494.96768, 488.6305, 479.9165, 470.88528, 461.616, 452.4255, 443.4723, 434.43948, 425.7232, 417.4028, 408.76508, 400.2855, 391.48856, 383.0875, 374.76538, 366.5222, 358.3579, 350.0348, 341.55276, 333.0704, 324.5877, 316.3425, 308.25552, 300.16824, 292.23923, 284.3892, 276.69748, 269.32266, 261.94757, 254.25499, 246.64145, 239.18623, 231.81007, 224.03705, 216.58102, 208.96606, 201.19218, 193.49734, 185.88153, 178.26546, 170.64908, 162.7944, 155.2568, 147.87762, 140.81558, 133.83264, 127.1669, 120.262856, 113.596664, 106.93026, 100.025536, 93.35869, 86.69162, 80.02434, 73.51559, 67.24477, 61.211903, 55.25824, 48.82809, 42.913765, 36.88018, 30.846416, 24.733082, 18.698963, 12.823464, 6.788993, 3.2158668, NaN, NaN, 499.08667, 494.4923, 488.55118, 480.07486, 470.64752, 461.29898, 452.4254, 443.63068, 435.07327, 426.4363, 417.8782, 409.31973, 400.84018, 392.51877, 384.11777, 376.03345, 367.94882, 359.78464, 351.6201, 343.37598, 335.29007, 327.3624, 319.35516, 311.50616, 303.4983, 295.4901, 287.4023, 279.31424, 271.2258, 263.13705, 254.9687, 246.40347, 238.07582, 230.0651, 222.13336, 214.20134, 206.42766, 198.65367, 190.87941, 183.2635, 175.568, 167.87218, 160.09674, 152.24167, 144.46564, 136.45125, 128.59526, 120.58027, 113.2792, 106.057236, 98.83502, 91.61255, 84.23108, 77.80184, 71.76929, 65.73656, 59.94179, 53.988094, 48.192993, 42.080177, 36.32444, 30.608232, 24.256706, 17.904984, 12.267663, 6.6301875, 2.1042144, NaN, NaN, 499.4033, 494.72974, 488.7886, 480.94604, 473.1032, 465.0224, 456.7828, 448.93906, 441.095, 433.1714, 425.16827, 417.24405, 409.3988, 401.39474, 393.6281, 386.099, 378.41104, 370.72284, 363.35138, 355.82114, 348.09244, 340.4031, 333.18912, 325.8956, 318.36398, 310.91138, 303.22064, 295.60892, 287.9969, 280.4639, 272.93063, 265.39706, 257.94254, 250.0912, 242.23958, 234.46695, 226.45609, 218.60355, 210.83003, 203.05623, 195.36145, 188.06305, 180.52638, 173.54482, 166.56299, 159.73962, 152.99538, 146.09221, 139.42686, 132.92, 126.65101, 119.90567, 113.39819, 106.89051, 100.144516, 93.557045, 87.36622, 81.01645, 74.90462, 69.18949, 63.752037, 58.35413, 53.03546, 47.875427, 42.556488, 36.99924, 31.600628, 25.963686, 20.326591, 14.848139, 8.813731, 3.2555664, NaN, NaN, 499.16534, 494.57098, 488.3922, 479.99512, 471.20157, 462.16998, 452.97952, 443.78867, 434.8351, 426.11887, 417.48154, 408.6853, 400.04724, 391.40878, 382.61148, 373.89304, 365.25348, 356.6136, 347.89404, 339.57053, 331.24664, 323.0017, 314.83572, 306.74872, 298.81995, 290.8116, 283.12012, 275.11115, 267.33978, 259.48883, 251.47893, 243.54805, 235.77548, 227.76466, 219.99152, 211.6628, 203.4924, 195.55966, 187.78528, 180.0106, 172.43398, 165.45212, 158.62872, 151.96379, 145.21928, 137.9191, 130.3806, 122.92118, 115.54085, 108.71578, 101.811134, 95.54118, 89.58853, 83.39758, 77.20645, 71.41202, 65.61742, 59.902035, 54.027725, 48.073864, 42.199215, 36.16562, 30.211235, 24.733051, 19.254719, 14.093839, 9.17103, 4.40691, 1.7071927, NaN, NaN, 501.26404, 496.74896, 490.88712, 482.807, 474.80582, 466.8835, 458.80246, 450.32495, 441.45093, 432.735, 424.0979, 415.46048, 406.90192, 397.86752, 389.0705, 380.11456, 371.15823, 362.2808, 353.3237, 344.52478, 335.5669, 326.60864, 317.72928, 309.32526, 301.00015, 292.51614, 284.19037, 275.94357, 268.09293, 260.47992, 252.9459, 245.64957, 238.0357, 230.5802, 223.28307, 215.50974, 207.57747, 199.56557, 191.55336, 183.46149, 175.36931, 166.95946, 159.10466, 151.09087, 143.07675, 135.06233, 127.68244, 120.461006, 113.47739, 106.65227, 99.66818, 93.001335, 86.41364, 79.666985, 73.39637, 67.20494, 60.77518, 54.424603, 48.15321, 42.119793, 36.32437, 31.163923, 25.52698, 19.572292, 13.935029, 9.012221, 4.3275037, 1.5483834, NaN, NaN, 498.6893, 493.61966, 487.124, 478.0139, 468.2696, 458.7625, 449.255, 440.064, 430.47638, 421.12604, 411.93378, 403.13736, 394.02353, 385.54337, 376.90433, 368.34418, 359.62515, 351.14355, 342.82016, 334.655, 326.37057, 317.9669, 309.56287, 301.39636, 293.46744, 285.1417, 276.97424, 268.64783, 260.63834, 252.5492, 244.8563, 237.1631, 229.8662, 222.48972, 215.50958, 208.44987, 201.38994, 194.25043, 187.34866, 180.04999, 172.9494, 165.88824, 159.06487, 152.24126, 145.41743, 138.83144, 132.40392, 125.8175, 119.151505, 112.4853, 106.29505, 100.18398, 94.31084, 88.5169, 82.80216, 77.16664, 71.68973, 66.371414, 60.814827, 55.09932, 49.423344, 43.945683, 38.547264, 33.70444, 28.9409, 24.733013, 19.889866, 14.967204, 11.156031, 7.5035896, 3.4540675, NaN, NaN, 499.75842, 495.1641, 488.90613, 480.03378, 470.44803, 461.17874, 452.3844, 443.51047, 434.79462, 425.52374, 416.88638, 408.4864, 399.61057, 390.57584, 381.937, 373.3771, 364.8168, 356.1769, 347.6952, 339.05457, 330.80997, 322.64432, 314.47833, 305.9949, 297.4318, 288.86838, 280.70105, 272.69202, 264.84125, 256.9902, 249.21817, 241.2872, 233.51457, 225.26573, 217.41318, 209.24303, 201.31052, 193.69504, 186.39659, 179.25656, 172.07661, 165.01543, 158.11267, 151.28905, 144.22714, 137.24434, 130.18196, 123.11933, 115.897736, 108.91397, 102.00934, 95.02511, 88.12, 81.37342, 74.86473, 68.35584, 62.00551, 56.13127, 50.177483, 44.382294, 38.66633, 33.18838, 27.789682, 22.787817, 17.706434, 12.863122, 8.257899, 3.3349612, NaN, NaN, 501.8968, 497.2233, 491.12384, 482.7269, 474.09192, 465.21893, 456.1871, 447.2341, 438.043, 429.16846, 420.2143, 411.10123, 401.9878, 393.34946, 384.71075, 376.0717, 366.8774, 358.55466, 350.4694, 342.3045, 334.06006, 325.57742, 317.1737, 308.76968, 299.96884, 291.40552, 283.3176, 275.07077, 266.9822, 258.89334, 250.96277, 243.11119, 235.41794, 227.88304, 220.34785, 212.89172, 205.356, 197.582, 190.12505, 182.42981, 174.6153, 166.91948, 159.14403, 151.36829, 143.43356, 135.49852, 127.959946, 120.50046, 113.8343, 106.92984, 100.18387, 93.834526, 87.32624, 80.897125, 74.467804, 68.11766, 61.687943, 55.019875, 48.748512, 43.112064, 37.991493, 32.98988, 28.226328, 23.70085, 19.413462, 14.887789, 9.171006, 3.6128697, NaN, NaN, 498.80707, 493.97507, 487.79633, 479.47845, 470.92258, 462.4456, 454.28516, 446.12442, 437.96335, 429.485, 421.24402, 413.16122, 405.0781, 396.91537, 388.67313, 380.50977, 372.26685, 364.1821, 356.09705, 348.2495, 340.52057, 332.75168, 325.14108, 316.89594, 308.72974, 300.95966, 293.34787, 285.8944, 278.51993, 271.14523, 263.77023, 255.99847, 248.54364, 241.08853, 233.3159, 225.38434, 217.61111, 209.59962, 201.8258, 194.21036, 186.51527, 179.05792, 171.6003, 163.98372, 156.92227, 149.86057, 142.87798, 136.21255, 129.46756, 123.19848, 117.008575, 110.9772, 105.26311, 99.46948, 93.834435, 88.04049, 82.32575, 76.45211, 70.73705, 64.94246, 59.147694, 53.194004, 47.875225, 43.112022, 38.904434, 34.696762, 30.409607, 25.884182, 22.152615, 17.54761, 12.148505, 5.95524, 2.0645027, NaN, NaN, 499.4799, 494.80637, 488.62762, 479.99292, 471.041, 462.0094, 452.97745, 443.78662, 434.83313, 425.95844, 417.24188, 408.2872, 399.17365, 390.29745, 381.8964, 373.3365, 364.77625, 356.37415, 347.97174, 339.56897, 331.16586, 322.2867, 313.24863, 305.0823, 296.6778, 287.95575, 279.07477, 270.11407, 261.54953, 253.06392, 244.41934, 236.17096, 228.08089, 220.22845, 212.2964, 203.65012, 195.32077, 187.38776, 179.1371, 170.8861, 162.91246, 154.9782, 147.12297, 139.42613, 131.49095, 124.03161, 117.04814, 110.54061, 104.11223, 97.52492, 90.54055, 83.55595, 76.5711, 69.9829, 63.473877, 57.04402, 50.613968, 44.183712, 38.1502, 32.910427, 27.749914, 22.43048, 17.825483, 13.220386, 7.8211718, 2.7394292, NaN, NaN, 499.51907, 494.6871, 488.42917, 479.8737, 471.31784, 462.524, 453.80896, 445.25204, 436.9325, 428.29562, 420.05463, 412.05103, 403.73013, 395.64664, 387.48358, 379.39948, 371.3943, 363.30954, 354.74887, 346.50494, 338.37958, 330.0557, 322.12787, 314.27905, 306.27133, 297.86688, 289.22418, 280.9776, 272.7307, 264.6421, 256.63245, 248.93973, 241.40533, 233.79137, 226.49437, 218.87984, 211.26503, 203.72926, 196.03456, 188.26024, 180.44595, 172.11569, 163.94376, 155.93019, 148.31303, 140.69562, 133.47467, 126.09475, 119.11136, 111.96901, 104.90578, 98.00103, 91.25479, 84.82582, 78.31727, 71.96726, 65.37892, 58.71099, 52.439762, 46.56527, 41.286022, 35.808167, 30.488945, 25.487164, 20.405865, 15.165642, 10.242887, 6.272836, 2.6997254, NaN, NaN, 499.95428, 495.12234, 488.8644, 480.62585, 472.86227, 464.62305, 456.3835, 448.0644, 439.74496, 431.34595, 423.10507, 414.86386, 406.30533, 398.22195, 390.21753, 382.45053, 374.68326, 366.99496, 359.4649, 351.85532, 344.40396, 337.1109, 329.65903, 321.8105, 314.27878, 307.06393, 299.4524, 291.91986, 284.38705, 276.69537, 269.00342, 261.46976, 254.01515, 246.56026, 239.18442, 232.04625, 224.7492, 217.53122, 210.07501, 202.8565, 195.4791, 188.10141, 180.5648, 172.86925, 165.25273, 157.79462, 150.2569, 143.03629, 135.65672, 128.67368, 122.08716, 115.65916, 109.5484, 102.80254, 96.29457, 90.10387, 84.23046, 78.03939, 71.37188, 64.38663, 57.83774, 51.725258, 46.406456, 41.246292, 36.086, 31.004967, 26.638355, 22.271648, 16.952082, 10.838378, 5.439111, 2.183602, NaN, NaN, 499.35965, 494.4485, 488.0321, 479.87274, 472.18835, 463.71146, 455.15497, 446.5189, 437.88245, 429.3249, 420.84622, 412.5257, 403.96707, 395.88364, 387.95834, 380.03278, 371.86914, 363.6259, 355.46158, 347.37622, 339.48874, 331.71985, 323.8714, 316.33975, 308.33215, 300.72067, 292.95032, 285.1797, 277.40875, 269.5582, 261.78668, 253.69765, 246.08414, 238.54967, 231.25285, 223.95578, 216.73778, 209.51952, 202.6183, 195.71686, 188.6962, 181.39761, 174.33678, 166.72034, 158.94492, 151.48659, 144.02798, 136.88652, 129.66545, 122.6822, 115.69871, 108.47689, 101.88974, 95.381744, 89.349754, 83.63508, 77.92024, 72.205246, 66.25196, 59.74283, 53.43195, 47.557503, 42.000435, 36.681385, 31.362198, 25.645903, 20.247032, 14.689222, 9.051862, 4.764188, 1.5880749, NaN, NaN, 499.00256, 494.01218, 487.67502, 479.67407, 472.14813, 463.98813, 456.0655, 447.7464, 439.58542, 431.3449, 423.34177, 415.2591, 407.01758, 399.0135, 391.40536, 383.5592, 375.71274, 367.94522, 360.25668, 352.4886, 344.68057, 337.07047, 329.46005, 321.84933, 314.39694, 306.6271, 299.09488, 291.40375, 283.71237, 276.09998, 268.88382, 261.42947, 253.89558, 246.91656, 239.85799, 232.56123, 225.26422, 217.72899, 210.35213, 202.81636, 195.24065, 187.46631, 179.85036, 172.3928, 164.69695, 157.23885, 150.09784, 142.87724, 135.81511, 128.99078, 122.40429, 115.97632, 109.78622, 103.6753, 97.64357, 91.61166, 85.18271, 78.991684, 72.64172, 66.92658, 61.1716, 55.218, 49.58176, 44.3423, 39.499653, 35.05384, 30.528542, 25.288595, 20.683683, 15.522883, 10.123754, 4.8832846, 1.6277745, NaN, NaN, 497.45743, 492.3878, 485.81293, 477.41583, 468.85992, 460.22443, 451.90552, 443.82394, 435.90054, 427.8976, 420.13208, 412.4455, 404.99637, 397.86395, 390.5728, 383.59845, 376.38605, 369.1734, 361.80197, 354.50955, 346.97906, 339.68613, 332.47217, 325.41656, 318.04355, 310.51175, 302.97964, 295.2887, 287.67673, 280.22308, 272.6106, 264.9978, 257.54333, 250.16792, 242.95085, 235.97147, 228.8332, 221.29813, 213.84207, 206.38576, 198.6912, 190.99632, 183.53918, 175.9231, 168.54474, 161.3248, 154.02527, 146.96352, 140.13956, 132.99797, 126.17356, 119.428276, 112.524055, 105.46087, 99.032364, 92.68303, 86.333496, 80.539375, 74.745094, 69.1094, 63.15603, 57.043728, 51.407547, 46.485683, 41.801865, 37.117943, 32.195736, 27.03523, 21.715805, 16.158049, 10.282542, 4.6450734, 1.6277728, NaN, NaN, 499.5165, 494.44693, 488.03058, 479.47513, 471.07776, 462.44238, 453.72742, 444.77438, 436.05865, 427.5803, 418.86386, 410.14703, 401.35062, 392.47455, 383.5981, 374.80057, 366.24042, 357.7592, 349.2776, 341.03345, 332.59082, 324.02893, 315.6252, 307.37976, 299.21326, 291.205, 283.27573, 275.18756, 267.17834, 259.32745, 251.63489, 244.02133, 236.4868, 228.87268, 221.3376, 213.72292, 206.10796, 198.41338, 190.79785, 183.26137, 176.12129, 168.90163, 161.6817, 154.30284, 146.60632, 138.83017, 130.73631, 122.80085, 115.02379, 107.40517, 100.103714, 93.04011, 86.37311, 80.023384, 73.67347, 67.24397, 61.052418, 55.336967, 49.541973, 43.826206, 38.665997, 33.108707, 27.233692, 21.596695, 16.435926, 12.069022, 6.193403, 2.2232943, NaN, NaN, 499.318, 494.40683, 488.0697, 479.1974, 470.16623, 461.21393, 452.41968, 443.54584, 434.75085, 426.0347, 417.3182, 408.44284, 399.5671, 390.8495, 382.21075, 373.3339, 365.01147, 356.68872, 348.36563, 339.72513, 331.441, 323.11688, 314.4753, 306.07123, 298.14255, 290.13428, 282.12567, 274.27536, 266.58334, 259.04965, 251.51567, 244.06075, 236.52621, 229.15005, 221.93227, 214.31761, 206.782, 199.08746, 191.23398, 183.38019, 175.68477, 167.75105, 160.21373, 152.99352, 145.93173, 138.79036, 131.49004, 124.03074, 116.967964, 109.825584, 102.60359, 95.46072, 88.555695, 81.57107, 74.66558, 67.99799, 62.044605, 56.01166, 50.296078, 44.580334, 38.94382, 33.862885, 28.62304, 22.906693, 17.348978, 12.346907, 7.900518, 3.533435, NaN, NaN, 499.47562, 494.88135, 488.9403, 480.781, 472.7006, 463.98608, 455.192, 446.4767, 437.7611, 429.12436, 420.408, 411.69128, 402.97418, 393.93973, 385.30112, 376.89996, 368.41916, 359.85876, 351.45657, 342.89548, 334.17548, 325.69293, 317.3686, 309.2025, 301.27396, 293.3451, 285.81238, 278.3587, 270.74615, 263.37125, 256.15466, 248.7792, 241.32417, 233.63094, 226.01674, 218.48157, 210.78748, 202.93445, 195.23978, 187.54482, 179.96857, 172.51105, 164.81523, 157.11914, 149.50209, 142.04346, 134.1878, 126.33185, 118.475586, 110.539665, 102.60343, 94.905, 87.60313, 80.380356, 73.31609, 66.330956, 59.90125, 53.630104, 47.914463, 42.51621, 36.998734, 32.076538, 26.519083, 20.564499, 14.689138, 9.76641, 4.6053567, 1.9056776, NaN, NaN, 500.4254, 495.75192, 489.73172, 481.01794, 471.9869, 463.3516, 454.9536, 446.79297, 438.7905, 430.6292, 422.15067, 413.751, 405.74722, 397.74316, 389.58026, 381.49628, 373.09497, 364.6933, 356.29132, 348.12677, 340.1601, 332.15347, 323.98798, 315.90143, 308.05243, 300.44098, 293.06714, 285.69302, 278.08075, 270.4682, 263.0933, 255.63878, 248.10472, 240.8083, 233.19437, 225.8181, 218.28294, 210.50954, 202.73582, 194.96184, 186.94955, 178.61961, 170.68604, 162.91083, 155.294, 147.43887, 139.90083, 132.44186, 124.90327, 117.443756, 110.14269, 102.92074, 95.698524, 88.63479, 81.49145, 74.66535, 68.31529, 62.20317, 56.170254, 50.137154, 44.540504, 38.66584, 32.71162, 26.67783, 21.279026, 16.356462, 11.910175, 5.6375694, 1.9850774, NaN, NaN, 498.16733, 493.25616, 486.8398, 478.36356, 469.9662, 461.48926, 452.85355, 444.21744, 435.34326, 427.1819, 418.94092, 410.62036, 402.458, 394.6123, 386.68704, 378.99927, 371.3112, 363.46432, 355.2208, 347.21478, 338.8517, 330.44867, 322.12454, 314.2758, 306.506, 298.73596, 290.64844, 282.87778, 275.424, 268.04926, 260.67426, 253.06108, 245.52692, 237.91318, 230.37846, 223.16074, 215.7048, 208.48657, 200.95078, 193.0974, 185.32304, 177.94507, 170.56683, 163.02965, 155.3335, 147.79576, 140.33708, 133.2749, 126.371185, 119.46724, 112.483696, 105.65864, 99.38891, 93.67456, 88.436264, 83.0391, 77.80053, 72.0062, 65.497314, 58.829453, 52.39953, 46.366325, 40.96805, 36.045963, 30.806196, 25.72508, 20.96142, 16.038857, 11.27497, 5.7963653, 2.1438801, NaN, NaN, 499.27576, 494.36462, 488.10675, 479.789, 471.62936, 463.15253, 454.59607, 446.11853, 437.71985, 429.08313, 420.68378, 412.2841, 403.88403, 395.24588, 386.7659, 378.3648, 369.88412, 361.08603, 352.4461, 343.96436, 335.72006, 327.7133, 319.86475, 311.85736, 303.84964, 295.8416, 287.754, 279.66605, 271.4985, 263.172, 255.00378, 247.07317, 239.22156, 231.21101, 223.75539, 216.53745, 208.76398, 201.06956, 193.29552, 185.8385, 178.38123, 171.003, 163.86255, 156.48381, 149.2635, 141.88425, 134.66342, 127.28363, 120.30036, 113.158134, 105.936295, 98.79357, 91.6506, 85.2217, 78.79261, 72.60145, 66.251335, 60.139168, 53.709286, 46.961666, 40.332905, 33.981792, 28.027447, 22.549295, 17.229792, 11.671953, 5.3993535, 1.9056704, NaN, NaN, 499.592, 494.7601, 488.58145, 480.0261, 471.2327, 462.2805, 453.16943, 444.2957, 435.9762, 427.41864, 419.25696, 410.6987, 402.4571, 394.21518, 386.1314, 378.1266, 370.12146, 361.87823, 354.1103, 346.57986, 339.04913, 331.5974, 324.14542, 316.77246, 309.55777, 302.10498, 294.9691, 287.59506, 280.2208, 272.68765, 265.07492, 257.6205, 250.32446, 242.86954, 235.57295, 228.1175, 220.74107, 213.36438, 205.82878, 198.29291, 190.47911, 182.46667, 174.1366, 166.04419, 157.95146, 150.1758, 142.39984, 134.70293, 126.926384, 119.546326, 112.483444, 105.6584, 98.67441, 91.84891, 85.10255, 78.75283, 72.641045, 66.529076, 60.337543, 54.14583, 47.834843, 41.56336, 35.60924, 29.813734, 24.494425, 19.49256, 14.887561, 9.567863, 4.1686263, 0.59552324, NaN, NaN, 499.35373, 494.28418, 487.70944, 478.8372, 469.8853, 460.53693, 451.02966, 441.52197, 432.25156, 422.9807, 413.78867, 404.04153, 394.69016, 385.17987, 376.0654, 366.6335, 357.5975, 348.3233, 338.89014, 330.01147, 321.25134, 312.4512, 303.9678, 295.80124, 287.71362, 279.54642, 271.45816, 263.0524, 255.0428, 247.19151, 239.49855, 231.8053, 224.03244, 216.10065, 208.08922, 200.39479, 192.54141, 184.52908, 176.43709, 168.5828, 160.80754, 153.032, 145.3355, 137.87677, 130.1797, 122.64106, 115.34022, 108.2772, 102.007576, 95.97585, 90.3408, 84.62621, 78.8321, 72.56158, 66.449615, 60.496227, 54.70143, 48.90647, 43.508278, 37.871777, 32.51299, 26.876186, 22.11257, 17.42824, 12.743802, 7.0270543, 2.739389, NaN, NaN, 499.98676, 495.39252, 489.29312, 480.97546, 472.57825, 464.02222, 455.22818, 446.35452, 437.79745, 429.0815, 420.20676, 411.41083, 402.6938, 393.89716, 385.2586, 376.54047, 368.05975, 359.2616, 350.78015, 342.37766, 334.45044, 326.44363, 318.59506, 310.98407, 303.2142, 295.60263, 287.8322, 279.98218, 271.97327, 264.04333, 256.03378, 248.26184, 240.80685, 233.82747, 227.00648, 220.50255, 213.6811, 206.62149, 199.32364, 191.78755, 184.44951, 177.30954, 170.328, 163.58424, 156.99895, 150.1754, 143.1136, 135.97218, 128.9099, 121.76799, 114.38777, 107.00728, 99.15034, 91.68993, 84.78485, 78.27639, 72.085236, 65.89388, 59.86111, 54.38383, 49.660553, 45.215015, 40.13428, 34.656475, 29.019741, 23.62103, 18.777948, 14.172946, 9.012043, 3.5334032, NaN, NaN, 500.22388, 495.23358, 488.73813, 479.78668, 470.99335, 461.64502, 452.21707, 442.78867, 433.59756, 424.80222, 416.00653, 407.36893, 398.81024, 390.09268, 381.61252, 373.132, 364.73038, 356.48697, 348.24323, 340.23697, 332.27005, 323.62894, 315.06677, 306.42496, 298.1792, 290.01242, 282.0832, 273.99506, 265.8273, 257.26273, 248.38055, 239.498, 231.01163, 222.68353, 214.75171, 206.89891, 199.04579, 191.19238, 183.81467, 176.43668, 169.49478, 162.35431, 155.37227, 148.46933, 141.64551, 134.90082, 128.23526, 121.56948, 114.74477, 108.078545, 101.6502, 95.14229, 89.03101, 83.55452, 78.07788, 72.12485, 65.77475, 59.6626, 53.550266, 47.358364, 41.245663, 35.529724, 29.972408, 24.891302, 20.048256, 14.8875065, 9.567828, 4.406815, 1.6277535, NaN, NaN, 499.23322, 494.55975, 488.61877, 480.85562, 473.80515, 466.2791, 458.83203, 451.4639, 444.25397, 436.5684, 428.72406, 420.8794, 412.95523, 405.26846, 397.42294, 389.49786, 381.81024, 373.726, 365.56226, 357.31888, 349.2337, 341.2275, 333.1417, 324.7385, 316.41418, 308.56528, 300.39893, 292.3908, 284.62027, 276.53223, 268.6025, 260.67245, 252.98003, 245.04938, 237.27704, 229.50441, 221.89012, 214.11693, 206.34341, 198.56963, 191.03352, 183.33847, 176.03981, 169.05824, 161.91776, 154.69768, 147.39801, 139.93938, 132.55981, 125.57677, 118.83156, 112.165474, 105.81663, 99.46758, 93.27708, 87.5626, 81.68922, 75.81567, 69.783195, 64.226814, 58.789356, 53.39144, 47.914, 41.9601, 36.482353, 30.925068, 25.129456, 19.651258, 14.093518, 9.250221, 4.4862113, 1.9453603, NaN, NaN, 501.094, 496.579, 490.40042, 481.9244, 473.52725, 464.49597, 455.4643, 446.353, 437.479, 428.44617, 419.33365, 410.0623, 401.1867, 392.70703, 384.06848, 375.4296, 366.55252, 357.27878, 348.32166, 339.20563, 330.00992, 320.97235, 312.09296, 303.0546, 294.49158, 286.16608, 277.84024, 269.27618, 261.18756, 253.25725, 245.40593, 237.63362, 229.86102, 222.00882, 214.31494, 206.54146, 198.60902, 190.75562, 182.74324, 174.49255, 166.43988, 158.10919, 149.77817, 141.28812, 133.2738, 125.89402, 118.8314, 111.92725, 105.102234, 98.594444, 91.92772, 85.498886, 78.9111, 72.95811, 67.08431, 61.607246, 56.130035, 50.25576, 43.984386, 38.18915, 32.949482, 27.947853, 23.025497, 17.467855, 11.274878, 4.6053066, 0.9528306, NaN, NaN, 498.3606, 493.37027, 486.95398, 478.87393, 471.26886, 463.42587, 455.18643, 447.10513, 439.0235, 431.10004, 422.93854, 414.856, 406.6146, 398.2144, 389.49683, 380.7789, 372.0606, 362.94565, 354.06808, 345.58646, 336.94595, 328.1465, 319.90167, 311.81506, 303.72815, 295.87875, 288.34622, 280.97205, 273.59756, 266.14352, 258.76852, 251.23465, 243.7798, 236.404, 229.02794, 221.49297, 213.79909, 205.78763, 197.77585, 189.44644, 181.4737, 173.46097, 165.84464, 158.228, 150.84912, 143.70802, 136.72537, 129.74248, 122.838715, 116.252144, 109.82407, 103.633896, 97.20544, 90.61804, 84.03043, 77.60136, 71.013336, 64.50447, 58.551064, 53.073776, 47.516956, 41.801216, 36.482258, 31.639502, 26.717241, 22.033043, 17.34874, 12.743726, 7.424011, 2.977577, NaN, NaN, 498.83536, 493.84506, 487.66644, 479.42798, 471.34763, 462.87085, 454.23526, 445.837, 437.35916, 428.80176, 420.244, 411.6066, 402.6519, 394.17227, 385.69232, 377.13275, 368.4143, 360.01257, 351.769, 343.68365, 335.91507, 327.74982, 319.6635, 311.73547, 303.80713, 296.03705, 288.66312, 280.89246, 272.96292, 265.42957, 258.05453, 250.44135, 242.43132, 234.26236, 226.01376, 217.92346, 210.15013, 202.21786, 194.68192, 187.14569, 179.68854, 172.07243, 164.21802, 156.12529, 148.11159, 140.49431, 132.9561, 125.65568, 118.593056, 111.76828, 105.57816, 99.62595, 93.51485, 87.32418, 81.92704, 76.13289, 70.2592, 64.70285, 59.46387, 54.14538, 48.70767, 42.674423, 36.402832, 30.607395, 25.28815, 20.206951, 15.205024, 9.726582, 4.3273935, 1.5483439, NaN, NaN, 501.25092, 496.5775, 490.399, 481.68533, 472.33755, 462.8309, 453.4823, 444.45016, 435.3384, 426.54318, 417.82684, 409.34787, 400.86853, 391.9926, 383.51257, 375.0322, 366.3929, 357.7533, 349.1926, 340.31442, 331.8719, 323.31012, 314.90652, 306.18546, 297.30545, 288.58362, 279.94073, 271.1389, 262.416, 254.0892, 246.00002, 238.30707, 230.53452, 222.52371, 214.75056, 206.8978, 198.41013, 190.1601, 182.06839, 174.0557, 166.51872, 159.29884, 152.2374, 145.41373, 138.11375, 130.73416, 122.719475, 115.101265, 108.038284, 101.37189, 94.70527, 88.117805, 81.53013, 74.86286, 68.59226, 62.242092, 56.44739, 50.652527, 44.698723, 38.903526, 32.869995, 27.153852, 21.675734, 16.118073, 10.639658, 5.2404976, 1.7468475, NaN, NaN, 500.4583, 495.7849, 489.76477, 482.08093, 474.55524, 466.55392, 458.39386, 449.9958, 441.59738, 433.43634, 425.1957, 416.63782, 408.3965, 400.31342, 392.38846, 384.701, 377.01324, 369.3252, 361.9539, 354.58234, 346.97275, 339.52136, 331.9112, 324.4593, 317.0864, 309.23755, 301.3091, 293.45966, 285.60992, 277.99774, 270.4646, 262.85187, 255.47676, 247.94278, 240.17061, 232.2395, 224.3081, 216.37639, 208.36505, 200.59137, 192.89673, 185.43977, 177.98257, 170.44576, 162.82932, 155.29193, 147.99232, 140.53375, 133.31296, 126.25061, 119.505455, 112.60136, 105.61767, 98.47501, 91.17337, 83.7921, 77.124916, 70.37814, 64.504295, 58.868427, 53.549923, 48.231285, 42.833122, 37.831757, 33.068436, 28.225613, 23.303284, 18.222044, 13.061281, 7.344592, 2.977569, NaN, NaN, 498.319, 493.64554, 487.70456, 480.17908, 472.4949, 464.57275, 456.6503, 448.72754, 440.96292, 433.1188, 425.43286, 417.6674, 410.13934, 402.69028, 395.08246, 387.7121, 380.3415, 372.9706, 365.59946, 357.91098, 350.61856, 343.24664, 335.71588, 328.50195, 321.1292, 313.67694, 306.22437, 299.00943, 291.7942, 284.42014, 277.04584, 269.59195, 262.2171, 254.9213, 247.38731, 239.93236, 232.31851, 224.46643, 216.61406, 208.76137, 201.06705, 193.53108, 186.07417, 178.93433, 171.79424, 164.8919, 158.06868, 151.0072, 144.50092, 137.91505, 131.40836, 125.139496, 118.94981, 112.998, 106.807945, 100.6177, 94.42727, 88.07791, 81.8871, 75.93423, 70.02086, 64.067635, 58.35238, 52.636963, 47.15954, 41.68197, 35.966087, 30.408827, 24.613237, 19.055668, 13.815536, 8.57527, 3.6524737, NaN, NaN, 498.87283, 494.041, 487.70395, 478.8318, 469.7216, 460.61096, 451.3415, 442.30933, 433.51443, 424.40222, 415.52734, 406.57285, 397.93494, 389.2174, 380.57877, 372.0983, 363.5382, 355.45334, 347.36816, 339.44122, 331.51398, 323.42786, 315.5, 307.88895, 300.51547, 292.98315, 285.4506, 278.3142, 270.93967, 263.72348, 256.34845, 249.13173, 241.51823, 233.82513, 226.68697, 219.70717, 212.48918, 205.35027, 197.97311, 190.35773, 182.74205, 174.88808, 167.27184, 159.73463, 152.35585, 144.9768, 137.59749, 130.29726, 123.39355, 116.4896, 109.58542, 102.76037, 95.69699, 89.34769, 83.31567, 77.28346, 71.33046, 65.37728, 59.26517, 53.073498, 47.15948, 41.443756, 35.96604, 30.805738, 25.724699, 20.405352, 15.16526, 9.925035, 4.684677, 1.7468412, NaN, NaN, 500.10013, 495.2683, 489.01056, 479.98, 471.02832, 462.0762, 453.20297, 444.40854, 435.9307, 427.611, 419.29092, 410.81204, 402.25357, 393.9325, 385.53183, 377.21005, 368.72946, 360.08997, 351.76718, 343.20627, 334.36752, 325.96442, 317.32315, 308.76077, 300.11877, 291.08, 282.19934, 273.23904, 264.43695, 255.63448, 246.91095, 238.34566, 229.46275, 221.13469, 213.04424, 204.95348, 197.10036, 189.40561, 181.55191, 173.6979, 165.68494, 157.67165, 149.49934, 141.16803, 132.91574, 124.58375, 116.64821, 108.95045, 101.56984, 94.82389, 88.395195, 82.12504, 75.93406, 70.13977, 64.504074, 58.86822, 53.152832, 47.754818, 42.197887, 37.117134, 32.115646, 26.87586, 21.238972, 15.998906, 10.520514, 5.3595743, 2.1835473, NaN, NaN, 500.575, 495.90164, 489.88153, 481.48477, 473.1669, 464.61102, 455.89633, 447.18127, 438.6243, 429.82928, 420.95465, 412.15887, 403.3627, 394.80392, 385.7693, 376.73425, 367.77805, 359.05927, 350.49866, 342.01697, 333.33673, 324.8543, 316.37155, 308.44342, 300.83212, 292.9827, 285.21225, 277.5208, 269.51187, 261.34402, 253.17587, 245.48323, 237.7903, 230.09708, 222.4829, 214.70978, 206.93637, 198.9247, 190.99203, 183.1384, 175.6018, 167.9856, 160.28976, 152.5143, 144.73853, 137.04182, 129.66223, 122.52045, 116.17198, 110.140755, 103.63319, 97.204765, 90.696785, 84.10922, 77.36271, 70.77472, 64.26589, 58.233143, 52.279594, 46.405254, 40.570442, 34.854546, 29.694223, 24.216202, 18.896824, 13.736099, 7.9400544, 3.017257, NaN, NaN, 499.06946, 494.2376, 487.8214, 478.87006, 469.36377, 459.93628, 451.14218, 442.5854, 434.02826, 425.3915, 416.59595, 407.95847, 399.47916, 391.39572, 383.23273, 375.22794, 367.30206, 358.97958, 350.73605, 342.1751, 333.81198, 325.3296, 316.76758, 308.2845, 299.95963, 291.55515, 283.3089, 274.98303, 266.5775, 258.33026, 250.00339, 241.8348, 234.22104, 226.60701, 219.15134, 211.93335, 204.55646, 196.70335, 189.2466, 181.94823, 174.72893, 167.58871, 160.36891, 153.30754, 145.92854, 138.31125, 131.01106, 123.86932, 116.965416, 110.29935, 103.633064, 97.12529, 91.014145, 85.22029, 79.66439, 73.87022, 67.996506, 62.122627, 56.248577, 50.453743, 44.777824, 39.220825, 33.425507, 27.709417, 22.548923, 17.467691, 12.54513, 7.1460543, 3.0966542, NaN, NaN, 498.94986, 494.19724, 488.1771, 480.09714, 472.17532, 463.93634, 455.53854, 447.3781, 439.45502, 431.05624, 422.81558, 414.81235, 406.6503, 398.4879, 390.4837, 382.16217, 374.15735, 366.15222, 357.90897, 349.74466, 341.6593, 333.49435, 325.1705, 317.0842, 308.99756, 301.22772, 293.37833, 285.6079, 277.83722, 270.7006, 263.56372, 256.5852, 249.44786, 242.31026, 235.41034, 228.19293, 221.45117, 214.47122, 207.25308, 199.95537, 192.73671, 184.88316, 177.26732, 169.6512, 162.11412, 154.89413, 147.91194, 141.0882, 133.78812, 126.963905, 120.377525, 114.029015, 107.36286, 100.775856, 94.268005, 88.077415, 82.04538, 76.33066, 70.695145, 65.05949, 59.542736, 53.986145, 48.429405, 42.872513, 37.236084, 31.917059, 26.677286, 21.357986, 16.435526, 11.512946, 5.716854, 2.1438391, NaN, NaN, 498.3551, 493.28564, 486.711, 477.83884, 468.6494, 459.61804, 450.03165, 440.99945, 432.2046, 423.1716, 413.97974, 405.10446, 396.30804, 387.5905, 378.79333, 370.47137, 362.3868, 354.6983, 346.61313, 338.28986, 330.28333, 322.5143, 314.50717, 306.6583, 298.8091, 290.72177, 283.03055, 274.94257, 267.2508, 259.8759, 252.42145, 244.88742, 236.87726, 229.34267, 222.04575, 214.9072, 207.7684, 200.86732, 193.64871, 186.42986, 178.8934, 171.35669, 163.42299, 155.489, 147.71338, 139.77878, 132.16125, 125.1783, 118.353806, 111.52908, 104.70414, 98.19642, 92.00596, 85.89468, 79.86259, 73.90969, 68.11537, 62.479645, 56.92314, 51.04896, 45.253998, 39.776413, 34.854404, 29.852882, 25.327593, 20.484629, 15.323965, 10.083775, 4.9228497, 1.6674302, NaN, NaN, 499.78046, 494.94864, 488.53247, 480.61102, 472.68924, 463.9749, 455.49792, 447.09982, 438.5429, 430.1441, 421.9034, 413.74167, 405.4211, 397.57568, 389.49222, 381.40845, 373.32434, 365.63623, 358.02707, 350.25912, 342.49088, 334.56378, 326.08148, 317.28168, 308.32297, 299.83957, 291.35583, 283.1096, 275.02164, 267.09195, 259.16196, 251.46959, 243.93553, 236.16327, 228.54933, 220.93513, 213.24132, 205.4679, 197.61485, 189.92017, 181.82854, 173.89525, 166.51703, 158.97986, 151.68044, 144.61879, 137.7156, 130.89154, 123.511765, 116.52851, 109.54501, 102.95809, 96.52969, 89.86298, 83.434166, 77.00515, 70.73468, 64.543396, 58.51068, 52.239643, 46.32564, 40.768707, 35.21162, 30.130722, 25.129091, 20.127338, 15.046067, 9.567679, 4.2479463, 1.5483271, NaN, NaN, 502.15625, 497.79977, 492.0174, 484.09604, 476.016, 467.46027, 458.74576, 449.8724, 440.8402, 431.41147, 421.98227, 412.6319, 402.80563, 393.1374, 383.70645, 374.51285, 365.3981, 356.3622, 347.48447, 338.84415, 330.3224, 321.8399, 313.43634, 305.03244, 296.7075, 288.69937, 280.61163, 272.52356, 264.4352, 256.1879, 248.01959, 240.00957, 232.31647, 224.46446, 216.8501, 208.83887, 200.82732, 192.9741, 184.96193, 177.02878, 169.13498, 161.43924, 153.7432, 146.36426, 139.2231, 132.24037, 125.01937, 117.95682, 111.21145, 104.62459, 98.59306, 92.40262, 85.97389, 79.78307, 73.75081, 67.639, 61.60638, 55.652966, 49.461227, 43.50746, 37.751987, 32.43299, 27.272638, 22.350334, 17.189728, 11.7908, 5.9947343, 2.1835327, NaN}
    CHLA = 
      {NaN, 0.138, 0.14100000000000001, 0.138, 0.138, 0.138, 0.138, 0.138, 0.14100000000000001, 0.11099999999999999, 0.138, 0.138, 0.135, 0.135, 0.11399999999999999, 0.132, 0.132, 0.135, 0.11699999999999999, 0.135, 0.138, 0.135, 0.135, 0.138, 0.10200000000000001, 0.132, 0.132, 0.135, 0.11099999999999999, 0.11099999999999999, 0.132, 0.135, 0.132, 0.11099999999999999, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.129, 0.135, 0.129, 0.132, 0.129, 0.135, 0.135, 0.135, 0.14400000000000002, 0.15300000000000002, 0.17400000000000002, 0.192, 0.237, 0.276, 0.324, 0.42900000000000005, 0.507, 0.723, 1.182, 1.02, 1.254, 0.363, 0.318, 0.30000000000000004, 0.28200000000000003, 0.237, 0.246, 0.237, NaN, NaN, 0.138, 0.138, 0.14100000000000001, 0.138, 0.138, 0.11699999999999999, 0.138, 0.138, 0.138, 0.138, 0.138, 0.138, 0.14100000000000001, 0.132, 0.129, 0.138, 0.135, 0.138, 0.135, 0.135, 0.10800000000000001, 0.135, 0.135, 0.135, 0.11099999999999999, 0.135, 0.10500000000000001, 0.135, 0.11099999999999999, 0.135, 0.135, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.129, 0.132, 0.132, 0.129, 0.129, 0.15000000000000002, 0.135, 0.14400000000000002, 0.15000000000000002, 0.17700000000000002, 0.195, 0.261, 0.30600000000000005, 0.339, 0.43499999999999994, 0.585, 0.735, 1.0470000000000002, 0.603, 0.30300000000000005, 0.273, 0.279, 0.261, 0.258, 0.24, NaN, NaN, 0.14400000000000002, 0.14100000000000001, 0.138, 0.135, 0.14100000000000001, 0.138, 0.138, 0.135, 0.135, 0.11399999999999999, 0.138, 0.135, 0.135, 0.129, 0.14100000000000001, 0.14100000000000001, 0.138, 0.11399999999999999, 0.14100000000000001, 0.135, 0.10800000000000001, 0.132, 0.135, 0.11099999999999999, 0.10800000000000001, 0.135, 0.135, 0.135, 0.11099999999999999, 0.132, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.129, 0.129, 0.11099999999999999, 0.129, 0.129, 0.11099999999999999, 0.10800000000000001, 0.132, 0.138, 0.14400000000000002, 0.15600000000000003, 0.165, 0.20700000000000002, 0.24, 0.237, 0.321, 0.35100000000000003, 0.43799999999999994, 0.684, 0.8699999999999999, 0.372, 0.23399999999999999, 0.29400000000000004, 0.246, 0.252, 0.23399999999999999, 0.22799999999999998, NaN, NaN, 0.138, 0.138, 0.138, 0.135, 0.14100000000000001, 0.14100000000000001, 0.135, 0.135, 0.132, 0.129, 0.138, 0.138, 0.135, 0.138, 0.132, 0.138, 0.132, 0.138, 0.135, 0.135, 0.135, 0.132, 0.135, 0.132, 0.132, 0.135, 0.11099999999999999, 0.132, 0.10800000000000001, 0.132, 0.132, 0.11099999999999999, 0.129, 0.129, 0.132, 0.132, 0.129, 0.10800000000000001, 0.10800000000000001, 0.129, 0.129, 0.135, 0.129, 0.129, 0.135, 0.129, 0.135, 0.129, 0.11099999999999999, 0.14100000000000001, 0.15300000000000002, 0.135, 0.20700000000000002, 0.279, 0.35700000000000004, 0.41100000000000003, 0.471, 0.603, 0.927, 0.42900000000000005, 0.264, 0.22799999999999998, 0.21600000000000003, 0.183, 0.21600000000000003, NaN, NaN, 0.138, 0.138, 0.135, 0.14100000000000001, 0.138, 0.138, 0.14100000000000001, 0.135, 0.135, 0.135, 0.126, 0.135, 0.11699999999999999, 0.138, 0.135, 0.135, 0.135, 0.135, 0.135, 0.132, 0.135, 0.132, 0.10500000000000001, 0.135, 0.135, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.10500000000000001, 0.129, 0.09, 0.132, 0.129, 0.10800000000000001, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.15300000000000002, 0.132, 0.132, 0.11099999999999999, 0.14100000000000001, 0.15600000000000003, 0.14400000000000002, 0.20700000000000002, 0.237, 0.321, 0.41700000000000004, 0.615, 0.96, 0.753, 0.381, 0.28800000000000003, 0.255, 0.23099999999999998, 0.23099999999999998, 0.24, 0.237, NaN, NaN, 0.138, 0.138, 0.135, 0.138, 0.14100000000000001, 0.14100000000000001, 0.135, 0.138, 0.138, 0.135, 0.138, 0.129, 0.138, 0.135, 0.14100000000000001, 0.135, 0.132, 0.132, 0.132, 0.132, 0.135, 0.135, 0.132, 0.138, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.11099999999999999, 0.129, 0.132, 0.129, 0.10500000000000001, 0.129, 0.10800000000000001, 0.129, 0.129, 0.10800000000000001, 0.129, 0.10800000000000001, 0.129, 0.132, 0.129, 0.129, 0.129, 0.10500000000000001, 0.132, 0.14100000000000001, 0.14400000000000002, 0.20400000000000001, 0.264, 0.33, 0.43200000000000005, 0.474, 0.744, 0.954, 0.96, 0.5760000000000001, 0.372, 0.30600000000000005, 0.258, 0.24, 0.198, 0.24, NaN, NaN, 0.138, 0.138, 0.138, 0.138, 0.11399999999999999, 0.135, 0.138, 0.138, 0.135, 0.132, 0.138, 0.126, 0.126, 0.10800000000000001, 0.138, 0.135, 0.132, 0.135, 0.135, 0.132, 0.138, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.135, 0.129, 0.132, 0.129, 0.129, 0.129, 0.129, 0.14100000000000001, 0.10800000000000001, 0.129, 0.132, 0.132, 0.11099999999999999, 0.129, 0.129, 0.10800000000000001, 0.11099999999999999, 0.14100000000000001, 0.168, 0.21000000000000002, 0.264, 0.333, 0.396, 0.5549999999999999, 0.726, 0.978, 0.684, 0.405, 0.22499999999999998, 0.237, 0.22199999999999998, 0.20400000000000001, 0.18, NaN, NaN, 0.14100000000000001, 0.138, 0.138, 0.14100000000000001, 0.138, 0.138, 0.138, 0.135, 0.09, 0.135, 0.132, 0.138, 0.11699999999999999, 0.138, 0.138, 0.138, 0.14100000000000001, 0.135, 0.138, 0.132, 0.135, 0.135, 0.135, 0.14100000000000001, 0.132, 0.135, 0.135, 0.132, 0.135, 0.11399999999999999, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.135, 0.132, 0.11099999999999999, 0.129, 0.132, 0.129, 0.132, 0.132, 0.129, 0.129, 0.129, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.135, 0.15000000000000002, 0.17700000000000002, 0.21300000000000002, 0.261, 0.35400000000000004, 0.498, 0.672, 0.792, 0.8160000000000001, 0.30600000000000005, 0.20400000000000001, 0.17400000000000002, 0.162, 0.15600000000000003, NaN, NaN, 0.138, 0.138, 0.138, 0.138, 0.138, 0.14100000000000001, 0.11099999999999999, 0.135, 0.138, 0.132, 0.132, 0.138, 0.138, 0.135, 0.138, 0.135, 0.10200000000000001, 0.10800000000000001, 0.135, 0.14100000000000001, 0.138, 0.135, 0.132, 0.135, 0.135, 0.11399999999999999, 0.135, 0.132, 0.135, 0.132, 0.135, 0.135, 0.135, 0.129, 0.129, 0.132, 0.11099999999999999, 0.132, 0.129, 0.132, 0.11099999999999999, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.129, 0.132, 0.11099999999999999, 0.135, 0.132, 0.132, 0.132, 0.138, 0.15300000000000002, 0.15600000000000003, 0.22499999999999998, 0.29100000000000004, 0.339, 0.42600000000000005, 0.5309999999999999, 0.627, 0.513, 1.149, 1.077, 0.795, 0.387, 0.267, 0.21300000000000002, 0.195, 0.171, 0.165, NaN, NaN, 0.135, 0.138, 0.138, 0.138, 0.138, 0.138, 0.135, 0.138, 0.135, 0.138, 0.135, 0.132, 0.11099999999999999, 0.11399999999999999, 0.138, 0.135, 0.135, 0.11399999999999999, 0.135, 0.135, 0.132, 0.135, 0.11399999999999999, 0.135, 0.135, 0.132, 0.132, 0.135, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.08700000000000001, 0.11099999999999999, 0.129, 0.129, 0.132, 0.129, 0.11099999999999999, 0.132, 0.15600000000000003, 0.132, 0.14100000000000001, 0.15600000000000003, 0.18, 0.23399999999999999, 0.28800000000000003, 0.33, 0.393, 0.387, 0.5549999999999999, 0.81, 1.119, 0.8640000000000001, 0.396, 0.324, 0.27, 0.28800000000000003, 0.186, NaN, NaN, 0.138, 0.135, 0.138, 0.14100000000000001, 0.138, 0.135, 0.135, 0.12, 0.132, 0.129, 0.129, 0.14100000000000001, 0.138, 0.138, 0.135, 0.135, 0.132, 0.135, 0.135, 0.132, 0.132, 0.132, 0.10500000000000001, 0.135, 0.132, 0.132, 0.10200000000000001, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.10800000000000001, 0.129, 0.129, 0.132, 0.126, 0.11099999999999999, 0.129, 0.129, 0.132, 0.129, 0.132, 0.132, 0.138, 0.14700000000000002, 0.159, 0.183, 0.22199999999999998, 0.261, 0.29400000000000004, 0.35100000000000003, 0.41700000000000004, 0.495, 0.675, 0.8550000000000001, 0.726, 0.42600000000000005, 0.44699999999999995, 0.33, 0.321, 0.31200000000000006, NaN, NaN, 0.138, 0.135, 0.135, 0.138, 0.138, 0.135, 0.138, 0.135, 0.129, 0.132, 0.11399999999999999, 0.126, 0.132, 0.138, 0.11699999999999999, 0.135, 0.081, 0.135, 0.135, 0.135, 0.138, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.129, 0.132, 0.129, 0.129, 0.132, 0.129, 0.10800000000000001, 0.129, 0.132, 0.10800000000000001, 0.11099999999999999, 0.129, 0.129, 0.129, 0.129, 0.132, 0.132, 0.132, 0.135, 0.14700000000000002, 0.162, 0.186, 0.23099999999999998, 0.27, 0.30000000000000004, 0.28800000000000003, 0.387, 0.43799999999999994, 0.5700000000000001, 0.642, 0.726, 0.43499999999999994, 0.43200000000000005, 0.396, 0.342, 0.264, 0.321, NaN, NaN, 0.135, 0.132, 0.135, 0.135, 0.135, 0.138, 0.138, 0.135, 0.135, 0.135, 0.126, 0.129, 0.11699999999999999, 0.135, 0.138, 0.138, 0.138, 0.135, 0.132, 0.132, 0.11099999999999999, 0.132, 0.135, 0.11099999999999999, 0.132, 0.135, 0.132, 0.135, 0.132, 0.132, 0.132, 0.10800000000000001, 0.11099999999999999, 0.132, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.10800000000000001, 0.132, 0.129, 0.129, 0.129, 0.132, 0.129, 0.132, 0.10800000000000001, 0.132, 0.14400000000000002, 0.135, 0.14400000000000002, 0.159, 0.171, 0.21000000000000002, 0.249, 0.30000000000000004, 0.30600000000000005, 0.43799999999999994, 0.558, 0.63, 0.8699999999999999, 0.519, 0.43499999999999994, 0.366, 0.315, 0.324, NaN, NaN, 0.135, 0.135, 0.132, 0.138, 0.135, 0.138, 0.132, 0.126, 0.126, 0.132, 0.132, 0.135, 0.135, 0.132, 0.138, 0.132, 0.135, 0.135, 0.11399999999999999, 0.135, 0.135, 0.135, 0.135, 0.10500000000000001, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.132, 0.132, 0.129, 0.132, 0.129, 0.132, 0.135, 0.14400000000000002, 0.15300000000000002, 0.159, 0.21899999999999997, 0.261, 0.28800000000000003, 0.255, 0.384, 0.51, 0.759, 0.759, 0.735, 0.44399999999999995, 0.366, 0.333, 0.315, 0.23399999999999999, NaN, NaN, 0.138, 0.138, 0.138, 0.138, 0.138, 0.11399999999999999, 0.138, 0.138, 0.11399999999999999, 0.135, 0.129, 0.126, 0.132, 0.132, 0.14100000000000001, 0.138, 0.135, 0.138, 0.10800000000000001, 0.135, 0.138, 0.138, 0.135, 0.135, 0.135, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.11099999999999999, 0.132, 0.129, 0.132, 0.129, 0.129, 0.129, 0.132, 0.132, 0.129, 0.129, 0.129, 0.132, 0.129, 0.132, 0.132, 0.132, 0.132, 0.14400000000000002, 0.165, 0.201, 0.21899999999999997, 0.273, 0.29100000000000004, 0.339, 0.387, 0.45899999999999996, 0.609, 0.741, 0.873, 0.43499999999999994, 0.35700000000000004, 0.29700000000000004, 0.30900000000000005, NaN, NaN, 0.138, 0.14100000000000001, 0.135, 0.135, 0.138, 0.135, 0.135, 0.132, 0.135, 0.138, 0.138, 0.135, 0.132, 0.129, 0.135, 0.138, 0.14100000000000001, 0.135, 0.135, 0.135, 0.135, 0.132, 0.135, 0.135, 0.135, 0.132, 0.132, 0.132, 0.135, 0.132, 0.132, 0.11099999999999999, 0.10800000000000001, 0.11099999999999999, 0.132, 0.132, 0.132, 0.129, 0.10500000000000001, 0.11099999999999999, 0.10800000000000001, 0.132, 0.129, 0.132, 0.129, 0.129, 0.126, 0.129, 0.129, 0.129, 0.129, 0.129, 0.132, 0.132, 0.14100000000000001, 0.15300000000000002, 0.17400000000000002, 0.20400000000000001, 0.249, 0.246, 0.276, 0.324, 0.31200000000000006, 0.396, 0.528, 0.768, 0.954, 1.332, 1.356, 0.636, 0.324, 0.28800000000000003, 0.22799999999999998, 0.246, NaN, NaN, 0.14100000000000001, 0.138, 0.135, 0.14100000000000001, 0.135, 0.135, 0.135, 0.138, 0.11399999999999999, 0.138, 0.138, 0.129, 0.14100000000000001, 0.138, 0.135, 0.138, 0.135, 0.138, 0.135, 0.135, 0.132, 0.132, 0.135, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.09, 0.132, 0.132, 0.129, 0.132, 0.10800000000000001, 0.129, 0.129, 0.129, 0.10800000000000001, 0.132, 0.10800000000000001, 0.129, 0.129, 0.132, 0.129, 0.138, 0.15000000000000002, 0.162, 0.189, 0.23399999999999999, 0.21600000000000003, 0.20700000000000002, 0.28200000000000003, 0.30600000000000005, 0.30900000000000005, 0.678, 0.8520000000000001, 1.332, 1.242, 0.9359999999999999, 0.396, 0.30600000000000005, 0.24, 0.21000000000000002, 0.21600000000000003, NaN, NaN, 0.132, 0.138, 0.138, 0.138, 0.138, 0.135, 0.138, 0.138, 0.138, 0.14100000000000001, 0.138, 0.11399999999999999, 0.129, 0.135, 0.135, 0.11099999999999999, 0.138, 0.135, 0.135, 0.135, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.10800000000000001, 0.132, 0.132, 0.129, 0.129, 0.10800000000000001, 0.129, 0.129, 0.129, 0.129, 0.132, 0.129, 0.10800000000000001, 0.132, 0.132, 0.138, 0.14400000000000002, 0.15300000000000002, 0.18, 0.237, 0.276, 0.28800000000000003, 0.327, 0.528, 0.687, 1.0050000000000001, 1.2480000000000002, 1.251, 1.287, 0.573, 0.30300000000000005, 0.261, 0.17700000000000002, 0.21899999999999997, NaN, NaN, 0.135, 0.135, 0.135, 0.132, 0.135, 0.135, 0.11399999999999999, 0.135, 0.138, 0.129, 0.14100000000000001, 0.135, 0.138, 0.135, 0.138, 0.135, 0.135, 0.135, 0.135, 0.135, 0.135, 0.135, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.10800000000000001, 0.132, 0.132, 0.132, 0.129, 0.129, 0.129, 0.132, 0.129, 0.132, 0.129, 0.129, 0.129, 0.129, 0.10500000000000001, 0.14100000000000001, 0.15000000000000002, 0.171, 0.198, 0.24, 0.279, 0.318, 0.393, 0.66, 0.867, 1.0350000000000001, 1.197, 1.221, 0.891, 0.35100000000000003, 0.30900000000000005, 0.28500000000000003, 0.261, NaN, NaN, 0.138, 0.135, 0.14100000000000001, 0.138, 0.135, 0.135, 0.138, 0.135, 0.135, 0.138, 0.11099999999999999, 0.129, 0.129, 0.14100000000000001, 0.135, 0.138, 0.138, 0.135, 0.135, 0.135, 0.11099999999999999, 0.135, 0.10800000000000001, 0.132, 0.135, 0.135, 0.132, 0.135, 0.132, 0.11399999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.11099999999999999, 0.132, 0.10800000000000001, 0.129, 0.10800000000000001, 0.135, 0.129, 0.129, 0.10800000000000001, 0.10800000000000001, 0.129, 0.129, 0.129, 0.129, 0.10800000000000001, 0.132, 0.11399999999999999, 0.14400000000000002, 0.129, 0.171, 0.189, 0.21300000000000002, 0.22499999999999998, 0.267, 0.327, 0.41700000000000004, 0.6990000000000001, 0.891, 1.131, 1.089, 0.5489999999999999, 0.42900000000000005, 0.339, 0.243, NaN, NaN, 0.138, 0.135, 0.135, 0.135, 0.135, 0.135, 0.135, 0.138, 0.135, 0.129, 0.138, 0.138, 0.138, 0.135, 0.138, 0.135, 0.135, 0.135, 0.132, 0.135, 0.132, 0.135, 0.135, 0.132, 0.11099999999999999, 0.132, 0.10500000000000001, 0.11099999999999999, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.132, 0.129, 0.129, 0.129, 0.129, 0.10500000000000001, 0.132, 0.132, 0.129, 0.11099999999999999, 0.138, 0.14700000000000002, 0.15300000000000002, 0.168, 0.183, 0.192, 0.22799999999999998, 0.249, 0.28500000000000003, 0.375, 0.489, 0.5820000000000001, 0.72, 0.783, 0.645, 0.489, 0.507, 0.396, 0.28800000000000003, 0.28500000000000003, NaN, NaN, 0.135, 0.135, 0.135, 0.135, 0.138, 0.135, 0.135, 0.132, 0.135, 0.135, 0.135, 0.129, 0.138, 0.132, 0.132, 0.138, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.135, 0.132, 0.132, 0.135, 0.132, 0.135, 0.132, 0.135, 0.132, 0.132, 0.129, 0.132, 0.10800000000000001, 0.132, 0.129, 0.129, 0.10800000000000001, 0.126, 0.129, 0.126, 0.10800000000000001, 0.129, 0.132, 0.129, 0.129, 0.132, 0.135, 0.12, 0.15300000000000002, 0.171, 0.189, 0.20700000000000002, 0.23099999999999998, 0.252, 0.30600000000000005, 0.366, 0.399, 0.498, 0.639, 0.756, 0.6900000000000001, 0.621, 0.399, 0.342, 0.243, 0.30300000000000005, NaN, NaN, 0.135, 0.132, 0.138, 0.138, 0.084, 0.11699999999999999, 0.135, 0.135, 0.135, 0.138, 0.10800000000000001, 0.132, 0.138, 0.132, 0.135, 0.135, 0.10800000000000001, 0.10800000000000001, 0.132, 0.135, 0.10800000000000001, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.11099999999999999, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.10800000000000001, 0.132, 0.129, 0.129, 0.129, 0.126, 0.129, 0.129, 0.129, 0.129, 0.132, 0.10500000000000001, 0.14100000000000001, 0.14700000000000002, 0.168, 0.17700000000000002, 0.17400000000000002, 0.21300000000000002, 0.237, 0.258, 0.29700000000000004, 0.40800000000000003, 0.5609999999999999, 0.666, 0.8370000000000001, 0.897, 0.8160000000000001, 0.5609999999999999, 0.43499999999999994, 0.399, 0.34500000000000003, NaN, NaN, 0.14100000000000001, 0.138, 0.11699999999999999, 0.138, 0.135, 0.14100000000000001, 0.11399999999999999, 0.138, 0.11099999999999999, 0.135, 0.135, 0.11099999999999999, 0.129, 0.132, 0.135, 0.138, 0.11399999999999999, 0.135, 0.132, 0.135, 0.135, 0.135, 0.132, 0.132, 0.11099999999999999, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.129, 0.10800000000000001, 0.129, 0.132, 0.129, 0.132, 0.129, 0.129, 0.126, 0.126, 0.129, 0.129, 0.138, 0.129, 0.129, 0.132, 0.138, 0.14700000000000002, 0.126, 0.14400000000000002, 0.195, 0.195, 0.20400000000000001, 0.21899999999999997, 0.21000000000000002, 0.31200000000000006, 0.45899999999999996, 0.6000000000000001, 1.242, 1.362, 0.8999999999999999, 0.75, 0.43200000000000005, 0.492, 0.44399999999999995, 0.498, 0.46199999999999997, NaN, NaN, 0.135, 0.138, 0.138, 0.138, 0.135, 0.135, 0.10800000000000001, 0.138, 0.135, 0.135, 0.11099999999999999, 0.135, 0.135, 0.132, 0.138, 0.135, 0.135, 0.132, 0.11099999999999999, 0.138, 0.132, 0.135, 0.132, 0.135, 0.135, 0.132, 0.132, 0.11099999999999999, 0.093, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.129, 0.126, 0.132, 0.132, 0.129, 0.129, 0.126, 0.129, 0.129, 0.129, 0.132, 0.138, 0.14400000000000002, 0.165, 0.17700000000000002, 0.183, 0.201, 0.23099999999999998, 0.21899999999999997, 0.46799999999999997, 0.567, 0.63, 0.7170000000000001, 0.897, 0.909, 1.059, 0.771, 0.471, 0.41700000000000004, 0.393, NaN, NaN, 0.138, 0.132, 0.138, 0.138, 0.132, 0.126, 0.126, 0.135, 0.138, 0.138, 0.138, 0.135, 0.135, 0.138, 0.132, 0.138, 0.135, 0.132, 0.135, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.129, 0.129, 0.132, 0.10800000000000001, 0.129, 0.129, 0.129, 0.129, 0.126, 0.10800000000000001, 0.129, 0.132, 0.126, 0.129, 0.129, 0.129, 0.129, 0.132, 0.132, 0.14700000000000002, 0.14400000000000002, 0.162, 0.17400000000000002, 0.189, 0.21300000000000002, 0.30000000000000004, 0.33, 0.6180000000000001, 0.639, 0.7080000000000001, 0.63, 0.5640000000000001, 1.002, 0.9510000000000001, 0.7110000000000001, 0.372, 0.28800000000000003, 0.24, 0.165, NaN, NaN, 0.135, 0.135, 0.138, 0.138, 0.138, 0.138, 0.132, 0.14100000000000001, 0.135, 0.129, 0.135, 0.14100000000000001, 0.135, 0.138, 0.135, 0.135, 0.135, 0.11099999999999999, 0.11099999999999999, 0.135, 0.11099999999999999, 0.132, 0.132, 0.11399999999999999, 0.135, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.129, 0.129, 0.11099999999999999, 0.126, 0.132, 0.10800000000000001, 0.129, 0.129, 0.129, 0.129, 0.132, 0.129, 0.132, 0.132, 0.138, 0.14100000000000001, 0.159, 0.17700000000000002, 0.186, 0.201, 0.21300000000000002, 0.28800000000000003, 0.43200000000000005, 0.45299999999999996, 0.46199999999999997, 0.684, 0.804, 0.6060000000000001, 0.762, 0.9119999999999999, 1.1099999999999999, 0.978, 0.396, 0.324, 0.27, 0.22799999999999998, NaN, NaN, 0.138, 0.132, 0.135, 0.138, 0.11699999999999999, 0.135, 0.135, 0.135, 0.135, 0.138, 0.132, 0.132, 0.138, 0.11099999999999999, 0.135, 0.132, 0.132, 0.10800000000000001, 0.135, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.10800000000000001, 0.10800000000000001, 0.11099999999999999, 0.132, 0.10800000000000001, 0.129, 0.129, 0.126, 0.129, 0.10500000000000001, 0.126, 0.129, 0.129, 0.10800000000000001, 0.132, 0.135, 0.159, 0.18, 0.189, 0.17700000000000002, 0.327, 0.399, 0.44099999999999995, 0.513, 0.492, 0.519, 0.6180000000000001, 0.774, 0.996, 1.056, 0.8520000000000001, 0.498, 0.42900000000000005, 0.405, 0.327, 0.35400000000000004, 0.003, NaN, NaN, 0.138, 0.14100000000000001, 0.138, 0.132, 0.10500000000000001, 0.135, 0.123, 0.132, 0.129, 0.138, 0.14100000000000001, 0.11399999999999999, 0.11099999999999999, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.11099999999999999, 0.132, 0.132, 0.11099999999999999, 0.132, 0.129, 0.129, 0.135, 0.129, 0.129, 0.126, 0.129, 0.129, 0.129, 0.129, 0.129, 0.135, 0.14400000000000002, 0.15300000000000002, 0.15600000000000003, 0.168, 0.168, 0.192, 0.273, 0.36, 0.46799999999999997, 0.477, 0.492, 0.474, 0.558, 0.651, 0.744, 0.75, 0.48, 0.30900000000000005, 0.381, 0.321, 0.315, 0.372, 0.43200000000000005, NaN, NaN, 0.135, 0.135, 0.135, 0.135, 0.135, 0.10800000000000001, 0.135, 0.138, 0.132, 0.129, 0.129, 0.10800000000000001, 0.11399999999999999, 0.135, 0.135, 0.11099999999999999, 0.132, 0.10800000000000001, 0.135, 0.132, 0.11099999999999999, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.10800000000000001, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.129, 0.132, 0.11099999999999999, 0.126, 0.129, 0.132, 0.135, 0.14100000000000001, 0.15000000000000002, 0.162, 0.15600000000000003, 0.168, 0.20400000000000001, 0.273, 0.336, 0.42600000000000005, 0.42900000000000005, 0.46499999999999997, 0.558, 0.627, 0.5489999999999999, 0.5760000000000001, 0.6060000000000001, 0.663, 0.513, 0.726, 0.534, 0.402, 0.384, 0.402, 0.321, 0.321, 0.387, NaN, NaN, 0.138, 0.135, 0.11099999999999999, 0.135, 0.135, 0.138, 0.132, 0.135, 0.135, 0.135, 0.129, 0.129, 0.10800000000000001, 0.135, 0.135, 0.132, 0.135, 0.132, 0.135, 0.132, 0.132, 0.10500000000000001, 0.135, 0.132, 0.11099999999999999, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.129, 0.132, 0.10800000000000001, 0.129, 0.135, 0.129, 0.129, 0.132, 0.10800000000000001, 0.10800000000000001, 0.132, 0.132, 0.138, 0.14400000000000002, 0.159, 0.18, 0.183, 0.20700000000000002, 0.264, 0.34500000000000003, 0.41100000000000003, 0.42600000000000005, 0.5609999999999999, 0.621, 0.609, 0.5640000000000001, 0.633, 0.5549999999999999, 0.657, 0.522, 0.378, 0.369, 0.369, 0.35700000000000004, 0.30900000000000005, NaN, NaN, 0.135, 0.138, 0.138, 0.135, 0.132, 0.135, 0.132, 0.132, 0.135, 0.126, 0.135, 0.132, 0.138, 0.135, 0.135, 0.138, 0.132, 0.135, 0.10800000000000001, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.129, 0.129, 0.129, 0.10800000000000001, 0.129, 0.129, 0.10800000000000001, 0.10800000000000001, 0.129, 0.129, 0.132, 0.135, 0.14100000000000001, 0.135, 0.18, 0.17700000000000002, 0.20700000000000002, 0.28200000000000003, 0.318, 0.384, 0.471, 0.5549999999999999, 0.552, 0.41100000000000003, 0.6000000000000001, 0.522, 0.645, 0.513, 0.513, 0.372, 0.35100000000000003, 0.29700000000000004, 0.35400000000000004, 0.36, 0.279, NaN, NaN, 0.135, 0.138, 0.135, 0.132, 0.129, 0.135, 0.135, 0.132, 0.135, 0.132, 0.138, 0.11399999999999999, 0.11699999999999999, 0.135, 0.132, 0.132, 0.135, 0.135, 0.11099999999999999, 0.132, 0.135, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.135, 0.135, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.129, 0.132, 0.129, 0.129, 0.10800000000000001, 0.10800000000000001, 0.135, 0.135, 0.138, 0.14700000000000002, 0.126, 0.168, 0.183, 0.21300000000000002, 0.29100000000000004, 0.36, 0.43499999999999994, 0.525, 0.5309999999999999, 0.54, 0.597, 0.642, 0.675, 0.579, 0.7050000000000001, 0.723, 0.5609999999999999, 0.489, 0.366, 0.36, 0.35400000000000004, 0.35400000000000004, 0.35700000000000004, 0.372, NaN, NaN, 0.138, 0.138, 0.10500000000000001, 0.135, 0.093, 0.138, 0.135, 0.135, 0.135, 0.132, 0.126, 0.132, 0.135, 0.135, 0.135, 0.11099999999999999, 0.135, 0.135, 0.135, 0.135, 0.138, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.132, 0.10800000000000001, 0.129, 0.132, 0.132, 0.129, 0.129, 0.132, 0.135, 0.135, 0.138, 0.15600000000000003, 0.162, 0.18, 0.18, 0.195, 0.261, 0.35100000000000003, 0.528, 0.579, 0.669, 0.6120000000000001, 0.522, 0.627, 0.6120000000000001, 0.627, 0.474, 0.318, 0.35400000000000004, 0.35100000000000003, 0.324, 0.30900000000000005, 0.28200000000000003, NaN, NaN, 0.135, 0.126, 0.126, 0.129, 0.126, 0.129, 0.132, 0.135, 0.138, 0.135, 0.132, 0.135, 0.10200000000000001, 0.138, 0.132, 0.135, 0.135, 0.132, 0.135, 0.132, 0.135, 0.132, 0.135, 0.11099999999999999, 0.132, 0.132, 0.132, 0.135, 0.132, 0.129, 0.132, 0.132, 0.10800000000000001, 0.11099999999999999, 0.132, 0.129, 0.129, 0.132, 0.132, 0.129, 0.129, 0.129, 0.132, 0.135, 0.138, 0.14100000000000001, 0.123, 0.15300000000000002, 0.168, 0.18, 0.186, 0.201, 0.22199999999999998, 0.255, 0.321, 0.375, 0.513, 0.5760000000000001, 0.6120000000000001, 0.678, 0.46799999999999997, 0.35400000000000004, 0.29100000000000004, 0.30000000000000004, 0.276, 0.237, 0.20400000000000001, 0.20400000000000001, 0.189, NaN, NaN, 0.135, 0.138, 0.138, 0.138, 0.11399999999999999, 0.135, 0.138, 0.135, 0.138, 0.138, 0.11399999999999999, 0.135, 0.135, 0.135, 0.135, 0.135, 0.132, 0.132, 0.11099999999999999, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.11399999999999999, 0.132, 0.135, 0.11099999999999999, 0.132, 0.132, 0.129, 0.129, 0.129, 0.132, 0.132, 0.10800000000000001, 0.11099999999999999, 0.129, 0.129, 0.129, 0.132, 0.132, 0.10800000000000001, 0.132, 0.132, 0.138, 0.14400000000000002, 0.14400000000000002, 0.15300000000000002, 0.162, 0.17400000000000002, 0.183, 0.20400000000000001, 0.22499999999999998, 0.249, 0.28200000000000003, 0.342, 0.43200000000000005, 0.46799999999999997, 0.534, 0.741, 0.492, 0.40800000000000003, 0.33, 0.342, 0.28500000000000003, 0.27, 0.252, 0.18, 0.195, 0.195, NaN, NaN, 0.138, 0.135, 0.135, 0.135, 0.138, 0.135, 0.135, 0.135, 0.11099999999999999, 0.129, 0.135, 0.135, 0.138, 0.135, 0.135, 0.135, 0.135, 0.135, 0.135, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.135, 0.129, 0.10800000000000001, 0.132, 0.129, 0.10800000000000001, 0.11399999999999999, 0.129, 0.132, 0.132, 0.135, 0.14400000000000002, 0.15000000000000002, 0.15600000000000003, 0.165, 0.18, 0.195, 0.22499999999999998, 0.20400000000000001, 0.279, 0.273, 0.46799999999999997, 0.43499999999999994, 0.627, 0.654, 0.78, 0.636, 0.43499999999999994, 0.399, 0.30600000000000005, 0.34500000000000003, 0.339, 0.30900000000000005, 0.23399999999999999, 0.246, NaN, NaN, 0.138, 0.126, 0.126, 0.129, 0.135, 0.132, 0.132, 0.138, 0.14100000000000001, 0.135, 0.135, 0.11399999999999999, 0.135, 0.11399999999999999, 0.135, 0.135, 0.135, 0.132, 0.132, 0.135, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.11399999999999999, 0.11099999999999999, 0.132, 0.132, 0.132, 0.129, 0.129, 0.129, 0.132, 0.129, 0.132, 0.10800000000000001, 0.132, 0.129, 0.132, 0.132, 0.132, 0.132, 0.132, 0.14100000000000001, 0.14400000000000002, 0.159, 0.171, 0.15600000000000003, 0.20400000000000001, 0.24, 0.28800000000000003, 0.34500000000000003, 0.381, 0.41400000000000003, 0.489, 0.6180000000000001, 0.687, 0.687, 0.5549999999999999, 0.34800000000000003, 0.36, 0.35100000000000003, 0.34500000000000003, 0.363, 0.35700000000000004, 0.39, 0.34500000000000003, NaN, NaN, 0.138, 0.135, 0.126, 0.126, 0.129, 0.129, 0.129, 0.138, 0.138, 0.11399999999999999, 0.135, 0.135, 0.10800000000000001, 0.135, 0.132, 0.132, 0.132, 0.135, 0.135, 0.135, 0.132, 0.11099999999999999, 0.132, 0.10800000000000001, 0.132, 0.132, 0.135, 0.132, 0.129, 0.132, 0.132, 0.132, 0.09, 0.132, 0.129, 0.129, 0.132, 0.11099999999999999, 0.129, 0.129, 0.129, 0.129, 0.10800000000000001, 0.129, 0.129, 0.129, 0.10800000000000001, 0.129, 0.129, 0.138, 0.138, 0.14700000000000002, 0.159, 0.171, 0.195, 0.20700000000000002, 0.255, 0.28200000000000003, 0.336, 0.43799999999999994, 0.495, 0.579, 0.7170000000000001, 0.675, 0.396, 0.34500000000000003, 0.372, 0.34800000000000003, 0.35100000000000003, 0.34500000000000003, 0.36, 0.342, 0.336, NaN, NaN, 0.132, 0.138, 0.135, 0.138, 0.138, 0.138, 0.138, 0.10800000000000001, 0.135, 0.135, 0.132, 0.135, 0.135, 0.135, 0.132, 0.135, 0.132, 0.135, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.129, 0.129, 0.132, 0.129, 0.129, 0.129, 0.129, 0.132, 0.11099999999999999, 0.129, 0.129, 0.10800000000000001, 0.10800000000000001, 0.129, 0.132, 0.129, 0.11099999999999999, 0.138, 0.12, 0.165, 0.171, 0.18, 0.189, 0.198, 0.22799999999999998, 0.243, 0.273, 0.336, 0.42600000000000005, 0.5309999999999999, 0.6060000000000001, 0.7020000000000001, 0.43799999999999994, 0.34800000000000003, 0.35700000000000004, 0.35400000000000004, 0.34500000000000003, 0.336, 0.336, 0.339, NaN, NaN, 0.138, 0.138, 0.138, 0.135, 0.135, 0.135, 0.135, 0.138, 0.135, 0.10800000000000001, 0.135, 0.132, 0.11099999999999999, 0.135, 0.132, 0.11399999999999999, 0.132, 0.135, 0.132, 0.132, 0.11099999999999999, 0.10500000000000001, 0.132, 0.10800000000000001, 0.132, 0.135, 0.132, 0.132, 0.129, 0.129, 0.129, 0.11099999999999999, 0.11099999999999999, 0.129, 0.129, 0.132, 0.129, 0.129, 0.132, 0.129, 0.129, 0.126, 0.129, 0.10800000000000001, 0.11099999999999999, 0.132, 0.14400000000000002, 0.15600000000000003, 0.165, 0.168, 0.17400000000000002, 0.15300000000000002, 0.201, 0.21899999999999997, 0.246, 0.279, 0.30900000000000005, 0.39, 0.534, 0.6120000000000001, 0.6240000000000001, 0.375, 0.342, 0.342, 0.35700000000000004, 0.339, 0.336, 0.342, NaN, NaN, 0.14100000000000001, 0.126, 0.129, 0.129, 0.132, 0.135, 0.11099999999999999, 0.135, 0.135, 0.135, 0.132, 0.135, 0.132, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.10800000000000001, 0.129, 0.129, 0.129, 0.129, 0.126, 0.129, 0.129, 0.10800000000000001, 0.129, 0.129, 0.10800000000000001, 0.132, 0.132, 0.132, 0.14100000000000001, 0.162, 0.165, 0.171, 0.192, 0.18, 0.24, 0.28500000000000003, 0.36, 0.43499999999999994, 0.579, 0.8699999999999999, 0.8490000000000001, 0.45299999999999996, 0.336, 0.33, 0.35400000000000004, 0.327, 0.27, 0.327, 0.339, NaN, NaN, 0.135, 0.132, 0.138, 0.135, 0.11399999999999999, 0.135, 0.132, 0.129, 0.138, 0.135, 0.135, 0.135, 0.132, 0.135, 0.135, 0.135, 0.132, 0.132, 0.132, 0.135, 0.11099999999999999, 0.11099999999999999, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.09, 0.132, 0.129, 0.129, 0.129, 0.132, 0.129, 0.132, 0.132, 0.132, 0.10800000000000001, 0.129, 0.129, 0.129, 0.129, 0.10500000000000001, 0.129, 0.129, 0.129, 0.129, 0.11099999999999999, 0.14100000000000001, 0.159, 0.165, 0.183, 0.20700000000000002, 0.249, 0.267, 0.29100000000000004, 0.387, 0.45899999999999996, 0.8370000000000001, 0.8999999999999999, 0.9750000000000001, 0.768, 0.43799999999999994, 0.30900000000000005, 0.30900000000000005, 0.30600000000000005, 0.21899999999999997, 0.246, NaN, NaN, 0.135, 0.132, 0.126, 0.135, 0.135, 0.135, 0.129, 0.138, 0.138, 0.138, 0.135, 0.10800000000000001, 0.11399999999999999, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.10800000000000001, 0.132, 0.11099999999999999, 0.129, 0.129, 0.132, 0.132, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.10800000000000001, 0.129, 0.129, 0.129, 0.10800000000000001, 0.129, 0.129, 0.10800000000000001, 0.135, 0.14100000000000001, 0.15600000000000003, 0.15600000000000003, 0.171, 0.186, 0.201, 0.186, 0.243, 0.258, 0.28200000000000003, 0.28200000000000003, 0.41700000000000004, 0.54, 0.8250000000000001, 0.7140000000000001, 0.8280000000000001, 0.678, 0.573, 0.258, 0.20700000000000002, 0.20700000000000002, 0.162, 0.192, NaN, NaN, 0.135, 0.135, 0.138, 0.135, 0.135, 0.132, 0.135, 0.138, 0.129, 0.135, 0.135, 0.135, 0.132, 0.135, 0.132, 0.135, 0.135, 0.132, 0.135, 0.132, 0.10800000000000001, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.129, 0.132, 0.129, 0.132, 0.129, 0.129, 0.132, 0.129, 0.129, 0.129, 0.129, 0.135, 0.126, 0.126, 0.129, 0.129, 0.129, 0.132, 0.132, 0.132, 0.135, 0.14400000000000002, 0.15600000000000003, 0.15600000000000003, 0.18, 0.186, 0.20700000000000002, 0.22199999999999998, 0.249, 0.28800000000000003, 0.36, 0.44999999999999996, 0.5820000000000001, 0.879, 0.996, 0.771, 0.399, 0.29400000000000004, 0.23399999999999999, 0.168, 0.195, NaN, NaN, 0.132, 0.129, 0.10500000000000001, 0.132, 0.132, 0.132, 0.129, 0.135, 0.138, 0.138, 0.135, 0.135, 0.135, 0.11399999999999999, 0.135, 0.132, 0.135, 0.135, 0.132, 0.10200000000000001, 0.132, 0.135, 0.132, 0.11099999999999999, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.132, 0.132, 0.129, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.135, 0.129, 0.129, 0.129, 0.132, 0.135, 0.135, 0.15000000000000002, 0.14700000000000002, 0.159, 0.17400000000000002, 0.186, 0.198, 0.22199999999999998, 0.24, 0.28200000000000003, 0.384, 0.507, 0.5309999999999999, 0.9630000000000001, 1.065, 1.0050000000000001, 0.675, 0.41100000000000003, 0.35700000000000004, 0.30900000000000005, 0.261, 0.237, NaN, NaN, 0.135, 0.132, 0.135, 0.138, 0.11099999999999999, 0.138, 0.135, 0.138, 0.135, 0.135, 0.11399999999999999, 0.135, 0.11399999999999999, 0.10800000000000001, 0.135, 0.132, 0.135, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.129, 0.129, 0.10800000000000001, 0.132, 0.129, 0.129, 0.129, 0.129, 0.10800000000000001, 0.129, 0.10800000000000001, 0.129, 0.132, 0.132, 0.11699999999999999, 0.14400000000000002, 0.14400000000000002, 0.162, 0.17700000000000002, 0.17700000000000002, 0.23099999999999998, 0.252, 0.30900000000000005, 0.31200000000000006, 0.399, 0.498, 0.732, 0.8190000000000001, 0.933, 0.8490000000000001, 0.5700000000000001, 0.474, 0.46799999999999997, 0.498, 0.489, 0.375, 0.48, NaN, NaN, 0.135, 0.135, 0.132, 0.132, 0.138, 0.138, 0.135, 0.132, 0.132, 0.132, 0.14100000000000001, 0.135, 0.135, 0.132, 0.135, 0.132, 0.135, 0.135, 0.132, 0.132, 0.11099999999999999, 0.11099999999999999, 0.132, 0.132, 0.10500000000000001, 0.09, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.10800000000000001, 0.129, 0.132, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.126, 0.129, 0.129, 0.132, 0.138, 0.14100000000000001, 0.14700000000000002, 0.15600000000000003, 0.165, 0.192, 0.21300000000000002, 0.22199999999999998, 0.24, 0.28200000000000003, 0.33, 0.399, 0.513, 0.7170000000000001, 0.9450000000000001, 0.654, 0.621, 0.384, 0.366, 0.369, 0.336, 0.378, 0.30300000000000005, NaN, NaN, 0.135, 0.132, 0.10500000000000001, 0.132, 0.135, 0.132, 0.135, 0.132, 0.132, 0.129, 0.11699999999999999, 0.138, 0.11399999999999999, 0.135, 0.132, 0.132, 0.135, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.10800000000000001, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.126, 0.132, 0.132, 0.10800000000000001, 0.132, 0.14100000000000001, 0.14700000000000002, 0.162, 0.17400000000000002, 0.186, 0.201, 0.20400000000000001, 0.21300000000000002, 0.22199999999999998, 0.249, 0.29100000000000004, 0.324, 0.369, 0.46799999999999997, 0.546, 0.66, 0.8759999999999999, 0.903, 0.591, 0.30000000000000004, 0.258, 0.31200000000000006, 0.30600000000000005, 0.29400000000000004, NaN, NaN, 0.132, 0.129, 0.132, 0.132, 0.10500000000000001, 0.123, 0.126, 0.129, 0.14100000000000001, 0.138, 0.10800000000000001, 0.135, 0.135, 0.135, 0.11099999999999999, 0.10800000000000001, 0.132, 0.132, 0.11099999999999999, 0.135, 0.132, 0.135, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.10800000000000001, 0.132, 0.11099999999999999, 0.132, 0.10800000000000001, 0.129, 0.129, 0.132, 0.10800000000000001, 0.126, 0.129, 0.10500000000000001, 0.126, 0.129, 0.135, 0.138, 0.14700000000000002, 0.14400000000000002, 0.129, 0.162, 0.183, 0.201, 0.21899999999999997, 0.246, 0.252, 0.28500000000000003, 0.34500000000000003, 0.43200000000000005, 0.522, 0.66, 0.8879999999999999, 0.642, 0.366, 0.318, 0.324, 0.318, 0.324, 0.44399999999999995, 0.402, 0.0, NaN, NaN, 0.34500000000000003, 0.333, 0.315, 0.321, 0.333, 0.327, 0.315, 0.30900000000000005, 0.31200000000000006, 0.318, 0.267, 0.318, 0.261, 0.30600000000000005, 0.30300000000000005, 0.31200000000000006, 0.30600000000000005, 0.264, 0.138, 0.135, 0.132, 0.11099999999999999, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.10800000000000001, 0.132, 0.129, 0.10800000000000001, 0.10800000000000001, 0.138, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.132, 0.132, 0.14400000000000002, 0.15600000000000003, 0.165, 0.17700000000000002, 0.192, 0.17700000000000002, 0.201, 0.267, 0.30000000000000004, 0.36, 0.44999999999999996, 0.5489999999999999, 0.7050000000000001, 0.759, 0.43799999999999994, 0.339, 0.35100000000000003, 0.30900000000000005, 0.315, 0.30300000000000005, 0.30600000000000005, 0.30600000000000005, NaN, NaN, 0.132, 0.135, 0.11099999999999999, 0.135, 0.132, 0.135, 0.138, 0.135, 0.10800000000000001, 0.132, 0.129, 0.129, 0.135, 0.135, 0.135, 0.135, 0.132, 0.135, 0.135, 0.132, 0.11099999999999999, 0.132, 0.10800000000000001, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.10800000000000001, 0.129, 0.132, 0.129, 0.132, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.10800000000000001, 0.132, 0.129, 0.11099999999999999, 0.129, 0.14400000000000002, 0.14400000000000002, 0.15300000000000002, 0.138, 0.186, 0.201, 0.22499999999999998, 0.243, 0.28500000000000003, 0.31200000000000006, 0.28500000000000003, 0.41100000000000003, 0.534, 0.879, 0.933, 0.795, 0.41100000000000003, 0.363, 0.321, 0.333, 0.29100000000000004, 0.29700000000000004, 0.273, NaN, NaN, 0.132, 0.138, 0.138, 0.138, 0.138, 0.138, 0.135, 0.138, 0.135, 0.132, 0.11399999999999999, 0.129, 0.135, 0.135, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.129, 0.126, 0.129, 0.129, 0.129, 0.129, 0.10800000000000001, 0.129, 0.129, 0.129, 0.129, 0.138, 0.14400000000000002, 0.15300000000000002, 0.138, 0.14700000000000002, 0.21000000000000002, 0.198, 0.261, 0.30300000000000005, 0.333, 0.363, 0.35700000000000004, 0.483, 0.567, 0.9119999999999999, 0.7050000000000001, 0.43200000000000005, 0.372, 0.35400000000000004, 0.252, 0.22799999999999998, 0.15300000000000002, 0.171, 0.159, NaN, NaN, 0.132, 0.132, 0.135, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.135, 0.135, 0.135, 0.135, 0.135, 0.132, 0.11099999999999999, 0.10500000000000001, 0.132, 0.132, 0.08700000000000001, 0.132, 0.132, 0.135, 0.11099999999999999, 0.129, 0.132, 0.132, 0.10800000000000001, 0.126, 0.132, 0.129, 0.132, 0.129, 0.129, 0.129, 0.129, 0.10800000000000001, 0.126, 0.129, 0.129, 0.129, 0.135, 0.14400000000000002, 0.15300000000000002, 0.165, 0.189, 0.22199999999999998, 0.249, 0.276, 0.30000000000000004, 0.35400000000000004, 0.327, 0.471, 0.651, 0.8400000000000001, 0.759, 0.46199999999999997, 0.363, 0.315, 0.27, 0.23399999999999999, 0.189, 0.183, 0.15600000000000003, NaN, NaN, 0.138, 0.135, 0.135, 0.135, 0.138, 0.10200000000000001, 0.11099999999999999, 0.132, 0.135, 0.135, 0.135, 0.11099999999999999, 0.132, 0.135, 0.132, 0.135, 0.138, 0.11099999999999999, 0.09, 0.132, 0.135, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.132, 0.129, 0.129, 0.129, 0.126, 0.126, 0.132, 0.129, 0.126, 0.126, 0.126, 0.132, 0.10800000000000001, 0.132, 0.138, 0.10800000000000001, 0.14700000000000002, 0.132, 0.171, 0.17700000000000002, 0.246, 0.258, 0.29100000000000004, 0.324, 0.30900000000000005, 0.42000000000000004, 0.585, 0.9870000000000001, 0.891, 0.483, 0.327, 0.30300000000000005, 0.29700000000000004, 0.261, 0.243, 0.249, 0.21899999999999997, NaN, NaN, 0.135, 0.135, 0.138, 0.135, 0.10500000000000001, 0.135, 0.138, 0.135, 0.132, 0.138, 0.132, 0.11399999999999999, 0.135, 0.132, 0.11099999999999999, 0.129, 0.135, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.10800000000000001, 0.132, 0.132, 0.129, 0.129, 0.132, 0.132, 0.132, 0.129, 0.129, 0.129, 0.129, 0.132, 0.132, 0.129, 0.126, 0.129, 0.10800000000000001, 0.10800000000000001, 0.10800000000000001, 0.129, 0.129, 0.10800000000000001, 0.129, 0.129, 0.129, 0.132, 0.138, 0.14700000000000002, 0.15600000000000003, 0.165, 0.171, 0.183, 0.198, 0.17700000000000002, 0.237, 0.246, 0.276, 0.342, 0.48, 0.5880000000000001, 0.8699999999999999, 1.008, 0.42000000000000004, 0.324, 0.30000000000000004, 0.28800000000000003, 0.23399999999999999, 0.27, NaN, NaN, 0.138, 0.135, 0.11099999999999999, 0.138, 0.135, 0.11099999999999999, 0.135, 0.135, 0.135, 0.11099999999999999, 0.132, 0.132, 0.132, 0.11099999999999999, 0.10200000000000001, 0.135, 0.135, 0.135, 0.135, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.129, 0.129, 0.132, 0.126, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.135, 0.135, 0.14400000000000002, 0.15300000000000002, 0.159, 0.171, 0.186, 0.189, 0.198, 0.22799999999999998, 0.246, 0.27, 0.29400000000000004, 0.41100000000000003, 0.528, 0.573, 0.879, 0.9690000000000001, 0.42300000000000004, 0.35700000000000004, 0.34500000000000003, 0.30300000000000005, 0.279, 0.267, 0.23099999999999998, NaN, NaN, 0.138, 0.135, 0.132, 0.135, 0.135, 0.138, 0.132, 0.132, 0.11099999999999999, 0.135, 0.09, 0.132, 0.132, 0.132, 0.132, 0.129, 0.11099999999999999, 0.135, 0.11099999999999999, 0.198, 0.135, 0.132, 0.135, 0.132, 0.11099999999999999, 0.099, 0.132, 0.132, 0.11099999999999999, 0.132, 0.129, 0.132, 0.10800000000000001, 0.129, 0.126, 0.132, 0.132, 0.126, 0.10800000000000001, 0.129, 0.129, 0.10800000000000001, 0.10800000000000001, 0.132, 0.135, 0.15000000000000002, 0.162, 0.135, 0.171, 0.195, 0.22799999999999998, 0.258, 0.28500000000000003, 0.34500000000000003, 0.46499999999999997, 0.552, 0.615, 0.8759999999999999, 0.801, 0.7050000000000001, 0.5369999999999999, 0.42300000000000004, 0.29700000000000004, 0.315, 0.273, 0.255, 0.129, NaN, NaN, 0.132, 0.138, 0.135, 0.138, 0.138, 0.135, 0.132, 0.132, 0.10800000000000001, 0.135, 0.132, 0.132, 0.138, 0.135, 0.126, 0.11399999999999999, 0.14100000000000001, 0.135, 0.132, 0.135, 0.135, 0.132, 0.132, 0.132, 0.11099999999999999, 0.11099999999999999, 0.11099999999999999, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.126, 0.10800000000000001, 0.129, 0.129, 0.132, 0.138, 0.12, 0.15600000000000003, 0.159, 0.138, 0.186, 0.201, 0.237, 0.252, 0.29400000000000004, 0.378, 0.477, 0.5940000000000001, 0.8310000000000001, 0.6990000000000001, 0.792, 0.579, 0.33, 0.327, 0.29400000000000004, 0.22499999999999998, 0.264, NaN, NaN, 0.135, 0.138, 0.135, 0.135, 0.138, 0.135, 0.138, 0.132, 0.10800000000000001, 0.135, 0.135, 0.132, 0.138, 0.135, 0.11399999999999999, 0.135, 0.132, 0.11099999999999999, 0.132, 0.135, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.129, 0.129, 0.129, 0.10800000000000001, 0.129, 0.10800000000000001, 0.129, 0.129, 0.129, 0.129, 0.129, 0.132, 0.132, 0.135, 0.123, 0.15300000000000002, 0.162, 0.168, 0.15600000000000003, 0.165, 0.21600000000000003, 0.23099999999999998, 0.255, 0.29700000000000004, 0.315, 0.387, 0.522, 0.753, 0.8130000000000001, 0.8759999999999999, 0.5940000000000001, 0.43200000000000005, 0.35100000000000003, 0.29700000000000004, 0.276, 0.28200000000000003, NaN, NaN, 0.135, 0.135, 0.135, 0.135, 0.132, 0.135, 0.135, 0.135, 0.138, 0.135, 0.135, 0.135, 0.11399999999999999, 0.11399999999999999, 0.129, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.132, 0.129, 0.129, 0.132, 0.129, 0.10800000000000001, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.10800000000000001, 0.129, 0.129, 0.10800000000000001, 0.132, 0.138, 0.14700000000000002, 0.159, 0.159, 0.17400000000000002, 0.195, 0.18, 0.22199999999999998, 0.237, 0.22199999999999998, 0.28500000000000003, 0.30900000000000005, 0.363, 0.471, 0.627, 0.765, 0.909, 0.729, 0.35100000000000003, 0.243, 0.273, 0.267, 0.28500000000000003, NaN, NaN, 0.135, 0.135, 0.135, 0.132, 0.132, 0.132, 0.11099999999999999, 0.135, 0.135, 0.132, 0.10500000000000001, 0.132, 0.132, 0.126, 0.11399999999999999, 0.138, 0.132, 0.135, 0.132, 0.132, 0.135, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.132, 0.129, 0.129, 0.129, 0.10800000000000001, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.129, 0.132, 0.14400000000000002, 0.15000000000000002, 0.159, 0.183, 0.20700000000000002, 0.22199999999999998, 0.22799999999999998, 0.24, 0.255, 0.28500000000000003, 0.321, 0.372, 0.43200000000000005, 0.63, 1.032, 0.762, 0.5760000000000001, 0.35400000000000004, 0.28200000000000003, 0.246, 0.252, 0.22199999999999998, 0.21600000000000003, NaN, NaN, 0.135, 0.135, 0.135, 0.138, 0.135, 0.135, 0.135, 0.132, 0.135, 0.135, 0.132, 0.09, 0.132, 0.135, 0.132, 0.11099999999999999, 0.129, 0.135, 0.138, 0.135, 0.135, 0.132, 0.135, 0.10500000000000001, 0.132, 0.132, 0.132, 0.132, 0.11099999999999999, 0.132, 0.132, 0.132, 0.132, 0.126, 0.129, 0.129, 0.126, 0.129, 0.129, 0.126, 0.129, 0.129, 0.132, 0.129, 0.129, 0.129, 0.129, 0.129, 0.135, 0.14400000000000002, 0.159, 0.168, 0.171, 0.17700000000000002, 0.23399999999999999, 0.27, 0.30300000000000005, 0.375, 0.48, 0.615, 0.909, 0.783, 0.5700000000000001, 0.44399999999999995, 0.375, 0.35700000000000004, 0.30600000000000005, 0.267, 0.23399999999999999, 0.0, NaN, NaN, 0.135, 0.132, 0.135, 0.138, 0.135, 0.135, 0.138, 0.135, 0.132, 0.10800000000000001, 0.11099999999999999, 0.135, 0.11399999999999999, 0.132, 0.132, 0.126, 0.132, 0.135, 0.10800000000000001, 0.135, 0.135, 0.10500000000000001, 0.132, 0.135, 0.11099999999999999, 0.132, 0.129, 0.132, 0.129, 0.132, 0.11099999999999999, 0.129, 0.11099999999999999, 0.10800000000000001, 0.129, 0.126, 0.129, 0.10800000000000001, 0.129, 0.126, 0.10800000000000001, 0.129, 0.126, 0.129, 0.135, 0.12, 0.15300000000000002, 0.162, 0.168, 0.14100000000000001, 0.18, 0.21000000000000002, 0.23099999999999998, 0.258, 0.31200000000000006, 0.372, 0.327, 0.525, 0.771, 0.759, 0.663, 0.489, 0.42900000000000005, 0.381, 0.321, 0.279, 0.258, 0.15600000000000003, NaN}
    DENSITY = 
      {NaN, 1029.1692, 1029.1427, 1029.1067, 1029.0624, 1029.0193, 1028.9786, 1028.9355, 1028.8921, 1028.8486, 1028.8048, 1028.7606, 1028.7152, 1028.666, 1028.6201, 1028.5745, 1028.5269, 1028.4758, 1028.4233, 1028.3743, 1028.3181, 1028.2625, 1028.201, 1028.1417, 1028.0828, 1028.0325, 1027.9742, 1027.925, 1027.8684, 1027.8033, 1027.7375, 1027.6691, 1027.6053, 1027.551, 1027.4867, 1027.4288, 1027.3672, 1027.3044, 1027.2437, 1027.1838, 1027.133, 1027.0844, 1027.0392, 1026.9934, 1026.9341, 1026.8678, 1026.8097, 1026.7512, 1026.6829, 1026.6034, 1026.499, 1026.4147, 1026.3171, 1026.1815, 1026.0497, 1025.908, 1025.7637, 1025.6163, 1025.4468, 1025.3005, 1025.21, 1025.0631, 1024.8735, 1024.6976, 1024.504, 1024.0001, 1023.8848, 1023.8632, 1023.8416, 1023.8107, 1023.7485, 1023.6697, NaN, NaN, 1029.1755, 1029.15, 1029.1144, 1029.0703, 1029.0214, 1028.973, 1028.923, 1028.8728, 1028.8184, 1028.7623, 1028.7045, 1028.6505, 1028.5973, 1028.5408, 1028.4891, 1028.4355, 1028.3871, 1028.337, 1028.2814, 1028.225, 1028.1692, 1028.1189, 1028.0659, 1028.0128, 1027.9519, 1027.89, 1027.8307, 1027.784, 1027.7233, 1027.647, 1027.5792, 1027.5167, 1027.4532, 1027.391, 1027.3378, 1027.2742, 1027.2101, 1027.1483, 1027.0984, 1027.0518, 1026.9996, 1026.9514, 1026.9044, 1026.8397, 1026.7753, 1026.702, 1026.6434, 1026.5668, 1026.4697, 1026.3052, 1026.1919, 1026.0151, 1025.7798, 1025.6061, 1025.4385, 1025.3528, 1025.2024, 1025.0825, 1024.9856, 1024.8121, 1024.252, 1023.89185, 1023.86487, 1023.83154, 1023.7938, 1023.7157, 1023.6681, NaN, NaN, 1029.1859, 1029.1592, 1029.1224, 1029.0802, 1029.0339, 1028.9915, 1028.949, 1028.9058, 1028.8591, 1028.8123, 1028.7609, 1028.7092, 1028.6583, 1028.6123, 1028.5659, 1028.5173, 1028.4664, 1028.4185, 1028.3583, 1028.3077, 1028.2651, 1028.2206, 1028.17, 1028.1119, 1028.0581, 1028.0109, 1027.9504, 1027.8881, 1027.8334, 1027.765, 1027.699, 1027.6313, 1027.5682, 1027.4991, 1027.4369, 1027.3773, 1027.3109, 1027.2369, 1027.1758, 1027.1171, 1027.0726, 1027.0251, 1026.975, 1026.916, 1026.8613, 1026.8015, 1026.7229, 1026.6752, 1026.636, 1026.5957, 1026.5002, 1026.3762, 1026.3038, 1026.1583, 1026.0826, 1025.9019, 1025.7396, 1025.5543, 1025.4001, 1025.2905, 1025.1554, 1024.9641, 1024.6863, 1023.94434, 1023.87823, 1023.795, 1023.7062, 1023.6709, 1023.6547, 1023.6381, NaN, NaN, 1029.163, 1029.1376, 1029.1025, 1029.051, 1029.0067, 1028.9601, 1028.9132, 1028.8599, 1028.8119, 1028.7528, 1028.6951, 1028.6426, 1028.5885, 1028.535, 1028.4845, 1028.43, 1028.3744, 1028.3175, 1028.267, 1028.2262, 1028.1759, 1028.1276, 1028.0834, 1028.0372, 1027.9893, 1027.929, 1027.8667, 1027.7933, 1027.7247, 1027.661, 1027.5695, 1027.4823, 1027.4067, 1027.3383, 1027.2671, 1027.2115, 1027.1583, 1027.1019, 1027.0377, 1026.9803, 1026.934, 1026.8827, 1026.8291, 1026.7761, 1026.7246, 1026.662, 1026.5891, 1026.5106, 1026.3997, 1026.3008, 1026.1891, 1026.0353, 1025.8595, 1025.6024, 1025.3729, 1025.2285, 1025.1212, 1025.0234, 1024.7526, 1024.269, 1023.81433, 1023.74274, 1023.71277, 1023.69086, 1023.67163, NaN, NaN, 1029.1683, 1029.1437, 1029.1108, 1029.0565, 1029.003, 1028.9496, 1028.8994, 1028.849, 1028.7982, 1028.7499, 1028.6964, 1028.6483, 1028.5973, 1028.5481, 1028.5051, 1028.4624, 1028.4188, 1028.3776, 1028.322, 1028.279, 1028.2318, 1028.1865, 1028.1423, 1028.0985, 1028.0514, 1028.0049, 1027.9569, 1027.8988, 1027.8243, 1027.744, 1027.6542, 1027.5494, 1027.4735, 1027.4015, 1027.3326, 1027.2783, 1027.2218, 1027.1649, 1027.1145, 1027.0677, 1027.0198, 1026.972, 1026.9165, 1026.8651, 1026.8134, 1026.7678, 1026.7201, 1026.6683, 1026.5908, 1026.5232, 1026.4346, 1026.3296, 1026.1858, 1026.0098, 1025.8589, 1025.7389, 1025.5248, 1025.2971, 1025.1311, 1024.8934, 1024.543, 1023.9742, 1023.85657, 1023.8282, 1023.73846, 1023.6863, 1023.65955, 1023.64105, NaN, NaN, 1029.1721, 1029.1488, 1029.114, 1029.0701, 1029.0253, 1028.977, 1028.9279, 1028.878, 1028.8307, 1028.7769, 1028.7256, 1028.677, 1028.6266, 1028.5831, 1028.536, 1028.4905, 1028.4456, 1028.4072, 1028.3666, 1028.3151, 1028.2695, 1028.226, 1028.1792, 1028.1417, 1028.0887, 1028.0375, 1027.9928, 1027.9406, 1027.8735, 1027.7782, 1027.667, 1027.5948, 1027.5266, 1027.4746, 1027.4222, 1027.3702, 1027.3029, 1027.2446, 1027.1945, 1027.15, 1027.1091, 1027.0659, 1027.0278, 1026.978, 1026.937, 1026.8953, 1026.8513, 1026.8102, 1026.7717, 1026.7278, 1026.6821, 1026.629, 1026.5845, 1026.5353, 1026.4379, 1026.2926, 1026.0813, 1025.912, 1025.6768, 1025.4646, 1025.2814, 1025.1235, 1024.9636, 1024.8044, 1024.519, 1024.12, 1023.86774, 1023.7276, 1023.60065, 1023.5649, 1023.54083, 1023.52203, NaN, NaN, 1029.1742, 1029.1505, 1029.1166, 1029.0676, 1029.0194, 1028.962, 1028.9154, 1028.871, 1028.8188, 1028.7745, 1028.7241, 1028.662, 1028.6089, 1028.5569, 1028.5087, 1028.4619, 1028.4156, 1028.3685, 1028.3201, 1028.2686, 1028.2264, 1028.1744, 1028.129, 1028.0747, 1028.0326, 1027.9917, 1027.9379, 1027.8829, 1027.8209, 1027.76, 1027.6779, 1027.5598, 1027.489, 1027.4337, 1027.3838, 1027.3414, 1027.269, 1027.2179, 1027.1671, 1027.1267, 1027.0851, 1027.0449, 1026.9929, 1026.9427, 1026.8966, 1026.8512, 1026.8053, 1026.7549, 1026.704, 1026.6519, 1026.6025, 1026.5474, 1026.4691, 1026.329, 1026.0933, 1025.8833, 1025.6525, 1025.4153, 1025.3103, 1025.1287, 1024.9828, 1024.8129, 1024.2734, 1023.83704, 1023.61743, 1023.5688, 1023.54614, 1023.5231, 1023.50714, NaN, NaN, 1029.1648, 1029.1348, 1029.0996, 1029.0538, 1029.0049, 1028.9613, 1028.9122, 1028.864, 1028.8148, 1028.7736, 1028.723, 1028.6732, 1028.6262, 1028.5723, 1028.525, 1028.4791, 1028.4307, 1028.384, 1028.3372, 1028.2931, 1028.2482, 1028.1901, 1028.148, 1028.1023, 1028.0541, 1028.003, 1027.9442, 1027.8807, 1027.814, 1027.7482, 1027.666, 1027.5975, 1027.5424, 1027.4861, 1027.4308, 1027.3789, 1027.3119, 1027.2556, 1027.2133, 1027.1674, 1027.1223, 1027.0774, 1027.028, 1026.9764, 1026.925, 1026.882, 1026.8364, 1026.7924, 1026.7496, 1026.701, 1026.6426, 1026.5897, 1026.5468, 1026.498, 1026.4164, 1026.2278, 1026.0156, 1025.8556, 1025.628, 1025.3663, 1025.1707, 1025.011, 1024.9296, 1024.6467, 1023.7673, 1023.5951, 1023.5674, 1023.54333, 1023.5276, NaN, NaN, 1029.146, 1029.1238, 1029.0875, 1029.0367, 1028.9856, 1028.9407, 1028.8993, 1028.8523, 1028.7997, 1028.7483, 1028.7006, 1028.6577, 1028.6112, 1028.5637, 1028.521, 1028.471, 1028.425, 1028.3773, 1028.3307, 1028.2863, 1028.243, 1028.1935, 1028.1478, 1028.0984, 1028.0482, 1027.9966, 1027.9401, 1027.8722, 1027.8071, 1027.7407, 1027.6652, 1027.5989, 1027.5339, 1027.4598, 1027.3969, 1027.3264, 1027.2645, 1027.2059, 1027.1509, 1027.104, 1027.057, 1027.0013, 1026.9565, 1026.917, 1026.8768, 1026.8422, 1026.8016, 1026.7587, 1026.7192, 1026.6721, 1026.605, 1026.5503, 1026.4908, 1026.3938, 1026.2357, 1026.053, 1025.8859, 1025.65, 1025.5145, 1025.3447, 1025.2389, 1025.1165, 1025.0729, 1024.8708, 1024.5765, 1024.281, 1023.96094, 1023.81287, 1023.6472, 1023.5995, 1023.5644, 1023.5474, NaN, NaN, 1029.1654, 1029.1412, 1029.1075, 1029.0558, 1029.0059, 1028.9562, 1028.908, 1028.8588, 1028.8114, 1028.7651, 1028.714, 1028.6647, 1028.6174, 1028.571, 1028.5256, 1028.4756, 1028.4263, 1028.3704, 1028.3151, 1028.2675, 1028.2129, 1028.1642, 1028.1136, 1028.0591, 1027.9991, 1027.9415, 1027.8746, 1027.8052, 1027.7184, 1027.6418, 1027.5693, 1027.4945, 1027.418, 1027.3344, 1027.2748, 1027.216, 1027.151, 1027.09, 1027.0358, 1026.9893, 1026.942, 1026.8947, 1026.8417, 1026.7924, 1026.739, 1026.6736, 1026.613, 1026.5469, 1026.4559, 1026.3419, 1026.1749, 1026.03, 1025.788, 1025.5862, 1025.4491, 1025.3019, 1025.1875, 1025.0931, 1024.924, 1024.6984, 1024.2584, 1023.9711, 1023.8839, 1023.746, 1023.6898, 1023.673, NaN, NaN, 1029.1487, 1029.1237, 1029.0916, 1029.0482, 1029.0065, 1028.9586, 1028.9078, 1028.8635, 1028.8131, 1028.7632, 1028.7177, 1028.6677, 1028.6174, 1028.5691, 1028.5211, 1028.476, 1028.4244, 1028.3649, 1028.316, 1028.2662, 1028.2103, 1028.1642, 1028.1113, 1028.0586, 1027.9922, 1027.932, 1027.8629, 1027.8007, 1027.7308, 1027.6606, 1027.5901, 1027.5309, 1027.4698, 1027.3993, 1027.3423, 1027.2777, 1027.2228, 1027.1724, 1027.1194, 1027.0667, 1027.0195, 1026.97, 1026.9215, 1026.8778, 1026.8204, 1026.7654, 1026.702, 1026.648, 1026.5826, 1026.5106, 1026.4059, 1026.2875, 1026.158, 1026.0055, 1025.8025, 1025.6444, 1025.5242, 1025.3441, 1025.1886, 1025.0754, 1024.9276, 1024.7799, 1024.5243, 1024.2762, 1024.0846, 1023.87024, 1023.8037, 1023.7901, NaN, NaN, 1029.1677, 1029.1434, 1029.1094, 1029.0646, 1029.0184, 1028.9723, 1028.9243, 1028.8759, 1028.8263, 1028.779, 1028.7303, 1028.6812, 1028.6338, 1028.5869, 1028.5371, 1028.4886, 1028.4376, 1028.3842, 1028.3301, 1028.2737, 1028.2211, 1028.1672, 1028.1158, 1028.0635, 1028.0054, 1027.945, 1027.8763, 1027.8087, 1027.7338, 1027.6709, 1027.5947, 1027.5294, 1027.4734, 1027.4104, 1027.3477, 1027.2937, 1027.2424, 1027.1902, 1027.1445, 1027.0999, 1027.0543, 1027.0094, 1026.9597, 1026.9102, 1026.8597, 1026.8097, 1026.7528, 1026.6895, 1026.626, 1026.5419, 1026.4299, 1026.3108, 1026.1776, 1026.0233, 1025.7766, 1025.6272, 1025.533, 1025.3938, 1025.2535, 1025.1377, 1025.0447, 1024.9355, 1024.744, 1024.3156, 1024.1367, 1024.0107, 1023.8475, 1023.80206, 1023.784, NaN, NaN, 1029.1576, 1029.1333, 1029.1023, 1029.0594, 1029.0208, 1028.9777, 1028.9354, 1028.8933, 1028.8527, 1028.8076, 1028.7603, 1028.7139, 1028.6683, 1028.6229, 1028.5775, 1028.5271, 1028.4778, 1028.4271, 1028.3739, 1028.3225, 1028.2661, 1028.2119, 1028.1595, 1028.108, 1028.0598, 1028.0023, 1027.9478, 1027.8921, 1027.8348, 1027.7657, 1027.7004, 1027.6505, 1027.6014, 1027.5435, 1027.4835, 1027.4241, 1027.3616, 1027.3156, 1027.2673, 1027.213, 1027.1635, 1027.1124, 1027.0652, 1027.0205, 1026.9783, 1026.9359, 1026.8853, 1026.8258, 1026.7687, 1026.706, 1026.6375, 1026.5531, 1026.4563, 1026.2983, 1026.1743, 1026.059, 1025.8602, 1025.6316, 1025.4669, 1025.2709, 1025.128, 1024.9955, 1024.8962, 1024.7458, 1024.4934, 1024.126, 1023.91504, 1023.81525, 1023.7751, NaN, NaN, 1029.145, 1029.1195, 1029.0857, 1029.0345, 1028.9829, 1028.9342, 1028.8871, 1028.8352, 1028.7844, 1028.7302, 1028.6758, 1028.623, 1028.5697, 1028.5166, 1028.4625, 1028.4126, 1028.3595, 1028.3021, 1028.2368, 1028.1843, 1028.1306, 1028.0801, 1028.0242, 1027.9714, 1027.9161, 1027.8605, 1027.8016, 1027.7487, 1027.6993, 1027.6406, 1027.5853, 1027.5325, 1027.4781, 1027.4261, 1027.3745, 1027.3235, 1027.2761, 1027.2295, 1027.1848, 1027.142, 1027.0912, 1027.0438, 1027.001, 1026.9556, 1026.9113, 1026.8514, 1026.7887, 1026.7283, 1026.6539, 1026.57, 1026.4425, 1026.3324, 1026.2253, 1026.0536, 1025.8256, 1025.6233, 1025.5044, 1025.3496, 1025.1732, 1025.0076, 1024.8411, 1024.6573, 1024.4689, 1024.2389, 1024.0206, 1023.9347, 1023.8607, 1023.8412, NaN, NaN, 1029.1492, 1029.1215, 1029.0884, 1029.0498, 1029.0139, 1028.9691, 1028.9237, 1028.8807, 1028.835, 1028.7948, 1028.755, 1028.712, 1028.6719, 1028.6276, 1028.5828, 1028.5383, 1028.4934, 1028.4467, 1028.4005, 1028.3567, 1028.308, 1028.2565, 1028.1981, 1028.1478, 1028.1024, 1028.0542, 1028.006, 1027.9518, 1027.9059, 1027.8431, 1027.7908, 1027.747, 1027.6931, 1027.6365, 1027.5867, 1027.5271, 1027.4681, 1027.4127, 1027.3625, 1027.3097, 1027.2576, 1027.2046, 1027.1523, 1027.1036, 1027.0526, 1027.0023, 1026.959, 1026.9082, 1026.8494, 1026.7993, 1026.7346, 1026.6631, 1026.5862, 1026.5011, 1026.4072, 1026.2792, 1026.1309, 1025.9117, 1025.7347, 1025.5848, 1025.4069, 1025.2306, 1025.124, 1025.0203, 1024.8887, 1024.7686, 1024.5468, 1024.1826, 1024.0707, 1023.9488, 1023.9311, NaN, NaN, 1029.1571, 1029.1313, 1029.0964, 1029.0533, 1029.0135, 1028.9673, 1028.9198, 1028.8761, 1028.832, 1028.7869, 1028.7405, 1028.6943, 1028.6447, 1028.6035, 1028.5591, 1028.5117, 1028.4639, 1028.4165, 1028.373, 1028.3282, 1028.2837, 1028.2301, 1028.1847, 1028.1362, 1028.0848, 1028.0294, 1027.9844, 1027.9243, 1027.8705, 1027.8135, 1027.76, 1027.6995, 1027.6418, 1027.5752, 1027.5234, 1027.4692, 1027.4022, 1027.3427, 1027.2941, 1027.2415, 1027.1915, 1027.1384, 1027.0939, 1027.0479, 1027.0007, 1026.9541, 1026.9015, 1026.8499, 1026.8031, 1026.7478, 1026.6853, 1026.6185, 1026.5297, 1026.4523, 1026.3247, 1026.167, 1026.0105, 1025.83, 1025.6753, 1025.5391, 1025.3936, 1025.2479, 1025.1235, 1025.0491, 1024.9805, 1024.847, 1024.7722, 1024.6646, 1024.5597, 1024.3468, 1023.939, 1023.78644, 1023.7678, 1023.7573, NaN, NaN, 1029.1614, 1029.135, 1029.1024, 1029.0491, 1028.9982, 1028.9484, 1028.8949, 1028.8455, 1028.7954, 1028.7422, 1028.6895, 1028.6354, 1028.5824, 1028.528, 1028.4634, 1028.4135, 1028.3545, 1028.298, 1028.2499, 1028.1941, 1028.1259, 1028.0717, 1028.0118, 1027.958, 1027.9019, 1027.8372, 1027.7782, 1027.7279, 1027.6727, 1027.6144, 1027.5461, 1027.4891, 1027.4243, 1027.3589, 1027.2935, 1027.2422, 1027.1833, 1027.1323, 1027.0769, 1027.0225, 1026.9767, 1026.9147, 1026.8618, 1026.814, 1026.7584, 1026.6906, 1026.597, 1026.4888, 1026.3759, 1026.265, 1026.129, 1025.9321, 1025.7273, 1025.5762, 1025.4703, 1025.3601, 1025.2689, 1025.0968, 1024.9313, 1024.7965, 1024.7043, 1024.6068, 1024.482, 1024.2108, 1023.9183, 1023.7907, 1023.7668, 1023.754, NaN, NaN, 1029.1713, 1029.147, 1029.1118, 1029.0625, 1029.0094, 1028.9603, 1028.9146, 1028.8674, 1028.8209, 1028.7697, 1028.7228, 1028.677, 1028.6288, 1028.5833, 1028.5267, 1028.4739, 1028.4172, 1028.3678, 1028.3137, 1028.2563, 1028.1962, 1028.1409, 1028.0807, 1028.0327, 1027.9756, 1027.916, 1027.8473, 1027.7753, 1027.7139, 1027.648, 1027.5851, 1027.5265, 1027.4767, 1027.4128, 1027.3552, 1027.305, 1027.2426, 1027.1869, 1027.1356, 1027.073, 1027.0172, 1026.959, 1026.8948, 1026.8282, 1026.7706, 1026.7084, 1026.6241, 1026.5254, 1026.4191, 1026.2972, 1026.1788, 1025.9957, 1025.7048, 1025.5209, 1025.3729, 1025.2651, 1025.0548, 1024.9423, 1024.8496, 1024.7288, 1024.6494, 1024.5686, 1024.3591, 1023.91486, 1023.7929, 1023.77, 1023.7468, NaN, NaN, 1029.1697, 1029.1454, 1029.1096, 1029.0603, 1029.0051, 1028.9531, 1028.905, 1028.856, 1028.8055, 1028.7571, 1028.7189, 1028.6675, 1028.616, 1028.564, 1028.5151, 1028.4567, 1028.4062, 1028.3563, 1028.304, 1028.249, 1028.196, 1028.1438, 1028.094, 1028.0448, 1027.9954, 1027.9386, 1027.8815, 1027.8319, 1027.7766, 1027.7173, 1027.6628, 1027.6069, 1027.5476, 1027.4888, 1027.4384, 1027.3906, 1027.334, 1027.2825, 1027.2281, 1027.1726, 1027.1234, 1027.0673, 1027.0106, 1026.9595, 1026.9054, 1026.8396, 1026.7694, 1026.7051, 1026.619, 1026.5236, 1026.4203, 1026.3141, 1026.2063, 1026.0543, 1025.8768, 1025.6666, 1025.4489, 1025.254, 1025.1088, 1024.951, 1024.8353, 1024.7734, 1024.687, 1024.6132, 1024.4962, 1023.932, 1023.79175, 1023.7573, 1023.732, NaN, NaN, 1029.1831, 1029.1561, 1029.1241, 1029.0797, 1029.0363, 1028.9889, 1028.9443, 1028.8949, 1028.8528, 1028.8044, 1028.7622, 1028.718, 1028.672, 1028.627, 1028.5809, 1028.5338, 1028.4866, 1028.4435, 1028.3958, 1028.3455, 1028.297, 1028.2471, 1028.2, 1028.1492, 1028.0977, 1028.0422, 1027.9929, 1027.9337, 1027.8881, 1027.838, 1027.7843, 1027.727, 1027.6832, 1027.6274, 1027.5667, 1027.5088, 1027.461, 1027.4053, 1027.3583, 1027.3016, 1027.2444, 1027.1921, 1027.1442, 1027.0979, 1027.0519, 1027.0077, 1026.9558, 1026.9021, 1026.8414, 1026.7856, 1026.7262, 1026.648, 1026.5708, 1026.465, 1026.3468, 1026.2434, 1026.1152, 1025.968, 1025.8467, 1025.6848, 1025.5466, 1025.3453, 1025.1854, 1025.0256, 1024.8217, 1024.7102, 1024.6442, 1024.5597, 1024.2833, 1023.9231, 1023.8376, 1023.7516, NaN, NaN, 1029.1763, 1029.1483, 1029.1118, 1029.061, 1029.0143, 1028.9644, 1028.9192, 1028.8701, 1028.82, 1028.7703, 1028.7213, 1028.674, 1028.6198, 1028.5724, 1028.5153, 1028.4598, 1028.4098, 1028.3596, 1028.3057, 1028.2474, 1028.188, 1028.1326, 1028.0762, 1028.0239, 1027.9667, 1027.9022, 1027.8359, 1027.7725, 1027.7152, 1027.652, 1027.5979, 1027.5345, 1027.4747, 1027.4159, 1027.3522, 1027.2826, 1027.2224, 1027.1661, 1027.0986, 1027.043, 1026.991, 1026.9401, 1026.8864, 1026.8257, 1026.7404, 1026.6538, 1026.5189, 1026.422, 1026.3168, 1026.1963, 1026.0472, 1025.8995, 1025.7365, 1025.5428, 1025.4354, 1025.2798, 1025.1069, 1024.9546, 1024.8342, 1024.7101, 1024.6062, 1024.3718, 1024.1425, 1024.0819, 1023.935, 1023.7736, 1023.75006, NaN, NaN, 1029.1794, 1029.1505, 1029.1177, 1029.0685, 1029.0231, 1028.9753, 1028.9269, 1028.8777, 1028.8314, 1028.7811, 1028.7352, 1028.6848, 1028.6368, 1028.5835, 1028.5269, 1028.4758, 1028.4305, 1028.3806, 1028.3301, 1028.2793, 1028.224, 1028.1677, 1028.1187, 1028.0638, 1028.0178, 1027.9642, 1027.9089, 1027.8516, 1027.7936, 1027.7311, 1027.6637, 1027.5996, 1027.5464, 1027.48, 1027.4172, 1027.3523, 1027.2905, 1027.235, 1027.174, 1027.1042, 1027.0413, 1026.9756, 1026.9144, 1026.8517, 1026.7819, 1026.7217, 1026.6476, 1026.5665, 1026.4463, 1026.2858, 1026.1469, 1025.9514, 1025.789, 1025.6614, 1025.5265, 1025.3491, 1025.1808, 1025.0754, 1025.0283, 1024.943, 1024.8013, 1024.6189, 1024.3984, 1024.1835, 1023.91547, 1023.8699, 1023.80664, 1023.7856, NaN, NaN, 1029.1896, 1029.1608, 1029.1215, 1029.0703, 1029.0181, 1028.9714, 1028.9177, 1028.8597, 1028.8134, 1028.7649, 1028.7109, 1028.6566, 1028.6062, 1028.5538, 1028.4993, 1028.4382, 1028.3795, 1028.3263, 1028.2668, 1028.206, 1028.1425, 1028.0911, 1028.032, 1027.9724, 1027.9215, 1027.8634, 1027.8081, 1027.7532, 1027.6991, 1027.6493, 1027.5859, 1027.5157, 1027.4583, 1027.3994, 1027.3402, 1027.2859, 1027.2235, 1027.1621, 1027.0916, 1027.0214, 1026.96, 1026.8967, 1026.8398, 1026.7751, 1026.7117, 1026.6469, 1026.5684, 1026.4885, 1026.3395, 1026.2008, 1026.0795, 1025.9396, 1025.8297, 1025.6188, 1025.3912, 1025.2867, 1025.1719, 1025.0354, 1024.9183, 1024.743, 1024.6052, 1024.4171, 1024.1296, 1023.9625, 1023.8959, 1023.85815, 1023.8325, NaN, NaN, 1029.1868, 1029.1573, 1029.1191, 1029.0673, 1029.0148, 1028.9662, 1028.9181, 1028.8702, 1028.8258, 1028.7709, 1028.7194, 1028.6669, 1028.6157, 1028.5686, 1028.5187, 1028.464, 1028.4082, 1028.3501, 1028.2916, 1028.2374, 1028.1774, 1028.1145, 1028.0629, 1028.0017, 1027.949, 1027.8955, 1027.8464, 1027.7914, 1027.7435, 1027.684, 1027.6309, 1027.5834, 1027.5309, 1027.4739, 1027.4047, 1027.3486, 1027.2817, 1027.2096, 1027.1366, 1027.0807, 1027.0215, 1026.9592, 1026.91, 1026.846, 1026.7761, 1026.707, 1026.6344, 1026.549, 1026.4702, 1026.3763, 1026.2361, 1026.068, 1025.9175, 1025.7474, 1025.6459, 1025.582, 1025.4459, 1025.3094, 1025.1434, 1025.0121, 1024.8901, 1024.7185, 1024.5698, 1024.4453, 1024.2147, 1023.9607, 1023.91345, 1023.8857, 1023.8691, 1023.85785, NaN, NaN, 1029.1975, 1029.1681, 1029.1279, 1029.0781, 1029.0214, 1028.9641, 1028.9106, 1028.8506, 1028.7933, 1028.7426, 1028.6963, 1028.6428, 1028.5966, 1028.5479, 1028.4976, 1028.4452, 1028.3904, 1028.3397, 1028.2864, 1028.2273, 1028.1759, 1028.1259, 1028.0714, 1028.0154, 1027.9613, 1027.8995, 1027.8439, 1027.7977, 1027.7428, 1027.6826, 1027.6237, 1027.5726, 1027.5187, 1027.4686, 1027.4185, 1027.3618, 1027.296, 1027.2314, 1027.1655, 1027.1138, 1027.0676, 1027.0013, 1026.9259, 1026.8491, 1026.777, 1026.7073, 1026.616, 1026.5508, 1026.4458, 1026.2981, 1026.1897, 1026.0323, 1025.882, 1025.7527, 1025.5916, 1025.3961, 1025.277, 1025.2002, 1025.1128, 1024.9832, 1024.8634, 1024.719, 1024.565, 1024.3972, 1024.0732, 1023.90753, 1023.8636, 1023.85504, NaN, NaN, 1029.1562, 1029.1302, 1029.092, 1029.0405, 1028.978, 1028.9205, 1028.863, 1028.8113, 1028.7606, 1028.7097, 1028.6593, 1028.607, 1028.5591, 1028.5066, 1028.4574, 1028.4082, 1028.3557, 1028.3035, 1028.2477, 1028.1958, 1028.141, 1028.0918, 1028.0381, 1027.9948, 1027.9481, 1027.8925, 1027.8348, 1027.7755, 1027.7155, 1027.6589, 1027.5941, 1027.5338, 1027.4674, 1027.4037, 1027.3438, 1027.2921, 1027.2316, 1027.1666, 1027.1033, 1027.0475, 1026.9763, 1026.9043, 1026.8237, 1026.7406, 1026.6462, 1026.5533, 1026.4719, 1026.3124, 1026.2006, 1026.0892, 1025.9348, 1025.7368, 1025.5707, 1025.4431, 1025.344, 1025.2213, 1025.1354, 1025.0767, 1024.9904, 1024.9012, 1024.8092, 1024.6816, 1024.2694, 1023.9551, 1023.9061, 1023.87744, 1023.85645, NaN, NaN, 1029.1758, 1029.1481, 1029.1133, 1029.0657, 1029.016, 1028.9684, 1028.9169, 1028.8668, 1028.8162, 1028.7618, 1028.7142, 1028.6687, 1028.6218, 1028.5748, 1028.5311, 1028.4807, 1028.4431, 1028.3931, 1028.3523, 1028.3019, 1028.2512, 1028.1951, 1028.152, 1028.1067, 1028.0614, 1028.0149, 1027.963, 1027.9095, 1027.854, 1027.8019, 1027.7494, 1027.694, 1027.6519, 1027.6078, 1027.5476, 1027.488, 1027.4271, 1027.3657, 1027.2979, 1027.244, 1027.1743, 1027.096, 1027.0326, 1026.9834, 1026.9174, 1026.8525, 1026.7694, 1026.6724, 1026.5773, 1026.5189, 1026.4073, 1026.2953, 1026.2002, 1026.012, 1025.8053, 1025.6649, 1025.567, 1025.4971, 1025.3615, 1025.2863, 1025.1816, 1025.1035, 1025.0612, 1024.9744, 1024.9038, 1024.8425, 1024.766, 1024.445, 1024.0774, 1023.9774, 1023.9327, 1023.9036, NaN, NaN, 1029.1805, 1029.1553, 1029.1173, 1029.069, 1029.0199, 1028.9607, 1028.9059, 1028.8479, 1028.791, 1028.7335, 1028.6744, 1028.6177, 1028.5646, 1028.5126, 1028.4591, 1028.4054, 1028.3455, 1028.2882, 1028.234, 1028.1793, 1028.1283, 1028.0758, 1028.0157, 1027.9574, 1027.8994, 1027.8347, 1027.787, 1027.7369, 1027.6823, 1027.6343, 1027.5793, 1027.5278, 1027.4651, 1027.3959, 1027.3438, 1027.2848, 1027.2097, 1027.1357, 1027.0872, 1027.0308, 1026.9509, 1026.8899, 1026.8169, 1026.7117, 1026.6201, 1026.5259, 1026.4625, 1026.3313, 1026.1969, 1025.9812, 1025.7748, 1025.6753, 1025.5076, 1025.418, 1025.3324, 1025.2681, 1025.1831, 1025.1208, 1025.0273, 1024.9358, 1024.8496, 1024.7957, 1024.6375, 1024.2732, 1024.1218, 1024.089, 1024.0626, 1024.0413, 1024.0255, NaN, NaN, 1029.1848, 1029.1586, 1029.1263, 1029.0797, 1029.033, 1028.9894, 1028.9386, 1028.8843, 1028.8232, 1028.7697, 1028.7166, 1028.6615, 1028.6094, 1028.5554, 1028.5059, 1028.4536, 1028.3972, 1028.339, 1028.2853, 1028.2313, 1028.1696, 1028.1077, 1028.0498, 1027.9966, 1027.9362, 1027.8861, 1027.8357, 1027.78, 1027.7263, 1027.6599, 1027.605, 1027.5557, 1027.4944, 1027.4288, 1027.3671, 1027.3079, 1027.2496, 1027.1743, 1027.0969, 1027.0222, 1026.9452, 1026.8601, 1026.797, 1026.6926, 1026.5703, 1026.455, 1026.3567, 1026.2714, 1026.1187, 1026.0065, 1025.7766, 1025.5859, 1025.4521, 1025.3501, 1025.2882, 1025.216, 1025.1306, 1025.0304, 1024.9199, 1024.7883, 1024.4597, 1024.2072, 1024.0574, 1024.0271, 1024.0, 1023.97797, 1023.9595, 1023.9478, NaN, NaN, 1029.1821, 1029.1494, 1029.114, 1029.0619, 1029.0035, 1028.951, 1028.893, 1028.8326, 1028.7716, 1028.7153, 1028.6611, 1028.6029, 1028.5459, 1028.4902, 1028.4369, 1028.3871, 1028.3323, 1028.2814, 1028.2322, 1028.1849, 1028.1299, 1028.0636, 1027.9972, 1027.9451, 1027.8967, 1027.8475, 1027.7969, 1027.7391, 1027.6813, 1027.6208, 1027.5647, 1027.5068, 1027.4462, 1027.3864, 1027.3365, 1027.2706, 1027.205, 1027.1428, 1027.0906, 1027.0243, 1026.9717, 1026.8892, 1026.8071, 1026.7275, 1026.6155, 1026.4857, 1026.3481, 1026.2236, 1026.1012, 1025.9678, 1025.7584, 1025.6193, 1025.5044, 1025.4159, 1025.3782, 1025.336, 1025.2253, 1025.1791, 1025.1307, 1025.0363, 1024.9379, 1024.8763, 1024.7485, 1024.4998, 1024.183, 1023.9789, 1023.9439, 1023.9219, 1023.9048, 1023.89136, 1023.87103, NaN, NaN, 1029.1858, 1029.1573, 1029.1213, 1029.0685, 1029.011, 1028.9476, 1028.895, 1028.8381, 1028.7864, 1028.7269, 1028.6664, 1028.6154, 1028.5627, 1028.5018, 1028.4465, 1028.3939, 1028.3472, 1028.2963, 1028.2389, 1028.18, 1028.1268, 1028.0781, 1028.029, 1027.9757, 1027.9241, 1027.8644, 1027.8102, 1027.7588, 1027.7083, 1027.6519, 1027.5975, 1027.5248, 1027.4562, 1027.397, 1027.3331, 1027.2743, 1027.205, 1027.1265, 1027.0599, 1026.9999, 1026.9211, 1026.8428, 1026.7756, 1026.6907, 1026.6147, 1026.5555, 1026.4056, 1026.2015, 1025.9674, 1025.8558, 1025.7576, 1025.6193, 1025.441, 1025.3905, 1025.335, 1025.2128, 1025.148, 1025.076, 1025.0066, 1024.9318, 1024.8145, 1024.4413, 1024.2046, 1023.99695, 1023.88434, 1023.8634, 1023.8428, 1023.82153, NaN, NaN, 1029.1948, 1029.166, 1029.1274, 1029.0748, 1029.0216, 1028.9712, 1028.9182, 1028.8636, 1028.8075, 1028.7511, 1028.6978, 1028.6467, 1028.5883, 1028.5283, 1028.4742, 1028.4222, 1028.3678, 1028.3112, 1028.2568, 1028.2, 1028.1472, 1028.0945, 1028.0369, 1027.9862, 1027.933, 1027.8815, 1027.8182, 1027.7584, 1027.7048, 1027.6467, 1027.5918, 1027.5367, 1027.4806, 1027.4279, 1027.364, 1027.2994, 1027.2196, 1027.1349, 1027.0757, 1027.0009, 1026.8961, 1026.8143, 1026.728, 1026.6462, 1026.5919, 1026.4554, 1026.2694, 1026.0674, 1025.9108, 1025.7495, 1025.5955, 1025.4999, 1025.4191, 1025.3711, 1025.2391, 1025.1768, 1025.0869, 1024.941, 1024.755, 1024.3647, 1024.2255, 1024.168, 1023.9261, 1023.8979, 1023.87946, 1023.8592, 1023.83356, 1023.8108, NaN, NaN, 1029.1675, 1029.1404, 1029.1057, 1029.0563, 1029.009, 1028.9551, 1028.9043, 1028.8574, 1028.8033, 1028.7555, 1028.7051, 1028.6572, 1028.6111, 1028.5543, 1028.5087, 1028.4622, 1028.4045, 1028.3447, 1028.2896, 1028.2406, 1028.1914, 1028.14, 1028.0898, 1028.0353, 1027.982, 1027.9286, 1027.8766, 1027.827, 1027.7761, 1027.7346, 1027.6748, 1027.6139, 1027.5706, 1027.5245, 1027.4678, 1027.4094, 1027.3501, 1027.294, 1027.2251, 1027.1544, 1027.0602, 1026.9844, 1026.9093, 1026.8153, 1026.7351, 1026.653, 1026.5546, 1026.458, 1026.3951, 1026.3022, 1026.1266, 1025.8882, 1025.7183, 1025.5677, 1025.4437, 1025.3804, 1025.2892, 1025.2438, 1025.2039, 1025.112, 1024.9886, 1024.8751, 1024.7819, 1024.5299, 1024.2328, 1024.1508, 1024.0128, 1023.9122, 1023.89624, 1023.8764, 1023.8522, 1023.82446, 1023.80707, NaN, NaN, 1029.1862, 1029.1577, 1029.1213, 1029.0662, 1029.0087, 1028.9565, 1028.903, 1028.8431, 1028.7948, 1028.7374, 1028.6874, 1028.6345, 1028.5844, 1028.5292, 1028.4723, 1028.4183, 1028.3611, 1028.3042, 1028.247, 1028.1869, 1028.1351, 1028.0839, 1028.0244, 1027.9806, 1027.9236, 1027.8613, 1027.8074, 1027.751, 1027.6958, 1027.633, 1027.5664, 1027.5089, 1027.4515, 1027.3881, 1027.3269, 1027.2561, 1027.1884, 1027.104, 1027.0259, 1026.897, 1026.817, 1026.7108, 1026.6183, 1026.5092, 1026.3898, 1026.241, 1026.0934, 1025.9578, 1025.7612, 1025.5919, 1025.451, 1025.2877, 1025.18, 1025.0975, 1024.9988, 1024.8987, 1024.7599, 1024.5753, 1024.2009, 1024.0054, 1023.9263, 1023.9017, 1023.8804, 1023.86084, 1023.8365, 1023.8162, NaN, NaN, 1029.1638, 1029.1355, 1029.0983, 1029.0469, 1028.9945, 1028.9388, 1028.8829, 1028.8317, 1028.7812, 1028.7324, 1028.6814, 1028.6278, 1028.5654, 1028.5167, 1028.4614, 1028.4126, 1028.3625, 1028.3141, 1028.2582, 1028.2034, 1028.1554, 1028.1055, 1028.0559, 1028.0011, 1027.953, 1027.9026, 1027.8441, 1027.7891, 1027.7338, 1027.6686, 1027.6138, 1027.5686, 1027.5195, 1027.4652, 1027.4034, 1027.34, 1027.2858, 1027.2297, 1027.1759, 1027.1055, 1027.041, 1026.939, 1026.8131, 1026.7075, 1026.6309, 1026.5183, 1026.4602, 1026.3019, 1026.1112, 1025.9744, 1025.8513, 1025.7029, 1025.5237, 1025.3385, 1025.1925, 1025.0951, 1024.9414, 1024.7386, 1024.4952, 1024.228, 1024.0293, 1023.96313, 1023.9395, 1023.9158, 1023.89435, 1023.86926, 1023.8471, 1023.82733, 1023.81024, NaN, NaN, 1029.1902, 1029.1611, 1029.1228, 1029.0737, 1029.0289, 1028.9749, 1028.9279, 1028.881, 1028.8293, 1028.777, 1028.7212, 1028.6656, 1028.614, 1028.5593, 1028.5105, 1028.457, 1028.4084, 1028.3527, 1028.3004, 1028.2468, 1028.1934, 1028.1489, 1028.1022, 1028.0461, 1027.9955, 1027.9426, 1027.8942, 1027.8438, 1027.7969, 1027.7421, 1027.6952, 1027.6469, 1027.6056, 1027.5464, 1027.4994, 1027.4542, 1027.3912, 1027.3367, 1027.2697, 1027.2057, 1027.1492, 1027.0782, 1027.0066, 1026.9103, 1026.7983, 1026.7008, 1026.6053, 1026.5238, 1026.4236, 1026.2891, 1026.1433, 1025.9758, 1025.837, 1025.6942, 1025.5471, 1025.4044, 1025.2699, 1025.164, 1025.0374, 1024.907, 1024.6117, 1024.3323, 1024.1156, 1024.0043, 1023.96454, 1023.94336, 1023.9226, 1023.905, 1023.88043, 1023.8523, 1023.8261, 1023.8115, NaN, NaN, 1029.1812, 1029.1514, 1029.1147, 1029.0685, 1029.0228, 1028.9728, 1028.9208, 1028.857, 1028.8026, 1028.7506, 1028.7006, 1028.6543, 1028.602, 1028.5466, 1028.4895, 1028.4403, 1028.3856, 1028.3297, 1028.271, 1028.2161, 1028.1682, 1028.1235, 1028.0723, 1028.0222, 1027.9695, 1027.9165, 1027.8705, 1027.8252, 1027.7776, 1027.723, 1027.6763, 1027.6271, 1027.5643, 1027.5114, 1027.4541, 1027.3896, 1027.3179, 1027.2499, 1027.2023, 1027.1411, 1027.0735, 1027.0027, 1026.9373, 1026.8657, 1026.7695, 1026.6735, 1026.6102, 1026.4425, 1026.3086, 1026.1672, 1026.0266, 1025.8534, 1025.6891, 1025.5658, 1025.4429, 1025.3059, 1025.1954, 1025.0071, 1024.8904, 1024.7971, 1024.5613, 1024.2981, 1024.1438, 1023.9922, 1023.95605, 1023.93176, 1023.9066, 1023.8817, 1023.8582, 1023.83905, 1023.82404, NaN, NaN, 1029.1747, 1029.1438, 1029.1088, 1029.0603, 1029.0145, 1028.9634, 1028.9164, 1028.868, 1028.8157, 1028.7656, 1028.7133, 1028.6611, 1028.6112, 1028.5619, 1028.5193, 1028.4694, 1028.4183, 1028.3661, 1028.3143, 1028.2539, 1028.2053, 1028.159, 1028.1135, 1028.0703, 1028.03, 1027.9797, 1027.9191, 1027.8667, 1027.8145, 1027.7594, 1027.7185, 1027.6609, 1027.6167, 1027.5625, 1027.4987, 1027.4375, 1027.3824, 1027.3098, 1027.2449, 1027.1903, 1027.1344, 1027.0798, 1027.011, 1026.9325, 1026.8448, 1026.7394, 1026.6619, 1026.5963, 1026.5177, 1026.4075, 1026.2728, 1026.112, 1025.9392, 1025.7723, 1025.6501, 1025.4929, 1025.3156, 1025.208, 1025.0868, 1024.9943, 1024.8965, 1024.762, 1024.5642, 1024.311, 1024.1206, 1023.96826, 1023.9488, 1023.92535, 1023.9047, 1023.8839, 1023.8574, 1023.83624, 1023.82166, NaN, NaN, 1029.1593, 1029.131, 1029.0953, 1029.0441, 1028.9888, 1028.9391, 1028.8876, 1028.8379, 1028.7869, 1028.7352, 1028.6838, 1028.632, 1028.583, 1028.5342, 1028.4878, 1028.4414, 1028.3905, 1028.3397, 1028.2959, 1028.2515, 1028.1969, 1028.1547, 1028.1086, 1028.0555, 1027.9983, 1027.9415, 1027.891, 1027.8416, 1027.7937, 1027.7428, 1027.695, 1027.6449, 1027.5884, 1027.5311, 1027.488, 1027.4336, 1027.378, 1027.3156, 1027.261, 1027.2025, 1027.1448, 1027.082, 1027.0139, 1026.9434, 1026.8927, 1026.836, 1026.7661, 1026.6956, 1026.6207, 1026.5261, 1026.4407, 1026.3022, 1026.0876, 1025.9001, 1025.7373, 1025.5935, 1025.3889, 1025.2887, 1025.1351, 1025.0038, 1024.8717, 1024.7676, 1024.5149, 1024.2118, 1024.0084, 1023.9721, 1023.9491, 1023.9285, 1023.9047, 1023.8798, 1023.8535, 1023.82825, 1023.81396, NaN, NaN, 1029.159, 1029.1261, 1029.0863, 1029.0332, 1028.9812, 1028.9276, 1028.8707, 1028.8193, 1028.7692, 1028.7108, 1028.6548, 1028.5975, 1028.5459, 1028.4878, 1028.4279, 1028.3812, 1028.3326, 1028.2819, 1028.2223, 1028.1613, 1028.0978, 1028.0361, 1027.9728, 1027.9193, 1027.863, 1027.8109, 1027.7559, 1027.6981, 1027.646, 1027.5868, 1027.5209, 1027.443, 1027.374, 1027.3215, 1027.2695, 1027.2142, 1027.151, 1027.0868, 1027.028, 1026.978, 1026.9215, 1026.8483, 1026.7742, 1026.7119, 1026.6234, 1026.5222, 1026.3927, 1026.1924, 1025.9541, 1025.8302, 1025.7118, 1025.6277, 1025.4678, 1025.3629, 1025.2731, 1025.1104, 1024.9867, 1024.8169, 1024.6573, 1024.3685, 1024.0446, 1023.9596, 1023.9318, 1023.90735, 1023.88513, 1023.86646, 1023.8388, 1023.8236, NaN, NaN, 1029.1371, 1029.111, 1029.077, 1029.024, 1028.968, 1028.9167, 1028.8645, 1028.7986, 1028.7456, 1028.6938, 1028.6426, 1028.5842, 1028.537, 1028.4727, 1028.4246, 1028.3707, 1028.3271, 1028.274, 1028.2163, 1028.1534, 1028.0953, 1028.0433, 1027.9822, 1027.9171, 1027.864, 1027.8121, 1027.7635, 1027.7141, 1027.6586, 1027.6044, 1027.5476, 1027.4843, 1027.4281, 1027.362, 1027.3007, 1027.2554, 1027.2091, 1027.1415, 1027.0764, 1027.0182, 1026.9629, 1026.901, 1026.8351, 1026.7534, 1026.6866, 1026.5782, 1026.4116, 1026.2687, 1026.1775, 1026.0608, 1025.8867, 1025.7188, 1025.6023, 1025.477, 1025.3478, 1025.2068, 1025.1117, 1025.0006, 1024.7893, 1024.591, 1024.3289, 1024.0027, 1023.9571, 1023.93225, 1023.9074, 1023.883, 1023.8678, 1023.84827, NaN, NaN, 1029.1714, 1029.1389, 1029.0961, 1029.038, 1028.9946, 1028.9481, 1028.8972, 1028.8398, 1028.7843, 1028.7279, 1028.6753, 1028.6188, 1028.5688, 1028.5161, 1028.4602, 1028.399, 1028.3503, 1028.2999, 1028.2451, 1028.1926, 1028.1333, 1028.0768, 1028.0215, 1027.9662, 1027.9114, 1027.8541, 1027.8055, 1027.7599, 1027.7108, 1027.6564, 1027.5988, 1027.5377, 1027.4756, 1027.415, 1027.3519, 1027.2893, 1027.2358, 1027.1799, 1027.122, 1027.0516, 1026.9823, 1026.9116, 1026.8466, 1026.7823, 1026.7211, 1026.6663, 1026.559, 1026.4015, 1026.2229, 1026.0459, 1025.8892, 1025.696, 1025.5189, 1025.3823, 1025.2083, 1025.0931, 1024.9626, 1024.823, 1024.6703, 1024.5255, 1024.208, 1024.0583, 1024.0374, 1024.0099, 1023.98517, 1023.9631, 1023.94086, 1023.9296, NaN, NaN, 1029.1836, 1029.1558, 1029.1136, 1029.0543, 1028.9955, 1028.948, 1028.9005, 1028.852, 1028.8014, 1028.7518, 1028.6954, 1028.6406, 1028.586, 1028.534, 1028.4664, 1028.4199, 1028.3743, 1028.3237, 1028.2745, 1028.2225, 1028.1666, 1028.1023, 1028.0475, 1027.9998, 1027.947, 1027.8889, 1027.8461, 1027.7942, 1027.7423, 1027.6909, 1027.6401, 1027.5775, 1027.5206, 1027.4705, 1027.4019, 1027.3458, 1027.2998, 1027.2382, 1027.167, 1027.1011, 1027.0297, 1026.9583, 1026.9003, 1026.8468, 1026.7988, 1026.7433, 1026.6813, 1026.6152, 1026.5299, 1026.3555, 1026.1882, 1025.9862, 1025.7817, 1025.5675, 1025.4209, 1025.2722, 1025.1736, 1025.0521, 1024.9094, 1024.7488, 1024.6533, 1024.5576, 1024.3197, 1024.1034, 1023.99316, 1023.9684, 1023.9484, 1023.92035, 1023.90393, NaN, NaN, 1029.1731, 1029.1462, 1029.102, 1029.048, 1028.9954, 1028.9409, 1028.8895, 1028.8362, 1028.7856, 1028.7313, 1028.6776, 1028.6267, 1028.5717, 1028.5138, 1028.4506, 1028.4033, 1028.3542, 1028.3015, 1028.2395, 1028.1805, 1028.1195, 1028.0634, 1028.0099, 1027.9557, 1027.907, 1027.8544, 1027.7999, 1027.7426, 1027.6887, 1027.6266, 1027.5808, 1027.5204, 1027.457, 1027.3997, 1027.361, 1027.316, 1027.2549, 1027.201, 1027.134, 1027.0681, 1027.0032, 1026.9427, 1026.8887, 1026.8381, 1026.7853, 1026.72, 1026.6536, 1026.543, 1026.3939, 1026.2443, 1026.0593, 1025.9247, 1025.764, 1025.6305, 1025.5178, 1025.3815, 1025.2657, 1025.1974, 1025.1222, 1024.9767, 1024.8376, 1024.7291, 1024.5986, 1024.4716, 1024.3936, 1024.2397, 1024.058, 1024.0283, 1023.99493, 1023.9702, 1023.9512, NaN, NaN, 1029.1759, 1029.1481, 1029.1128, 1029.0605, 1029.0045, 1028.9513, 1028.8955, 1028.8472, 1028.8046, 1028.7516, 1028.702, 1028.655, 1028.5936, 1028.5371, 1028.4747, 1028.4054, 1028.3513, 1028.2933, 1028.2341, 1028.1885, 1028.14, 1028.0881, 1028.0325, 1027.9769, 1027.9141, 1027.8588, 1027.8036, 1027.7511, 1027.7013, 1027.6426, 1027.5856, 1027.5264, 1027.4674, 1027.3998, 1027.3419, 1027.2906, 1027.2299, 1027.16, 1027.0939, 1027.0283, 1026.9617, 1026.907, 1026.8556, 1026.802, 1026.7432, 1026.6777, 1026.606, 1026.4799, 1026.339, 1026.2015, 1026.036, 1025.8806, 1025.7302, 1025.5747, 1025.4062, 1025.285, 1025.1787, 1025.0883, 1024.9268, 1024.7795, 1024.6182, 1024.503, 1024.4182, 1024.1951, 1024.0236, 1023.9866, 1023.95844, 1023.9405, NaN, NaN, 1029.1825, 1029.1509, 1029.1149, 1029.0629, 1029.0045, 1028.9451, 1028.8911, 1028.8317, 1028.7743, 1028.7228, 1028.6632, 1028.6147, 1028.5698, 1028.516, 1028.462, 1028.407, 1028.3542, 1028.3053, 1028.2546, 1028.2087, 1028.1611, 1028.114, 1028.0559, 1028.0021, 1027.9531, 1027.896, 1027.8439, 1027.7886, 1027.7347, 1027.6877, 1027.6387, 1027.5874, 1027.5267, 1027.4637, 1027.4005, 1027.3584, 1027.3154, 1027.267, 1027.1973, 1027.1217, 1027.0497, 1026.995, 1026.9349, 1026.867, 1026.8046, 1026.7401, 1026.656, 1026.5741, 1026.4542, 1026.3015, 1026.1902, 1026.0219, 1025.8519, 1025.7457, 1025.6329, 1025.5048, 1025.3184, 1025.178, 1025.043, 1024.9073, 1024.7993, 1024.6747, 1024.5739, 1024.441, 1024.2689, 1024.0455, 1024.0138, 1023.99066, 1023.9644, 1023.94684, NaN, NaN, 1029.1604, 1029.1326, 1029.091, 1029.0378, 1028.9882, 1028.9314, 1028.8657, 1028.8058, 1028.7484, 1028.6954, 1028.6383, 1028.5835, 1028.5239, 1028.4645, 1028.4062, 1028.3402, 1028.2755, 1028.212, 1028.1564, 1028.1079, 1028.061, 1028.0132, 1027.9498, 1027.8937, 1027.8376, 1027.781, 1027.7216, 1027.6532, 1027.5986, 1027.5339, 1027.4624, 1027.4008, 1027.3386, 1027.2798, 1027.2336, 1027.1729, 1027.1019, 1027.0233, 1026.9672, 1026.8888, 1026.8345, 1026.7563, 1026.6697, 1026.5709, 1026.4443, 1026.3246, 1026.1753, 1026.0184, 1025.879, 1025.6669, 1025.4832, 1025.3357, 1025.2207, 1025.1044, 1025.0023, 1024.9131, 1024.7571, 1024.6635, 1024.5411, 1024.4181, 1024.1974, 1024.0804, 1024.0559, 1024.035, 1024.0161, 1023.98987, 1023.97064, NaN, NaN, 1029.188, 1029.1615, 1029.123, 1029.0707, 1029.0215, 1028.9698, 1028.918, 1028.8657, 1028.814, 1028.7615, 1028.7047, 1028.6465, 1028.5948, 1028.5375, 1028.4801, 1028.4236, 1028.3668, 1028.3108, 1028.253, 1028.1915, 1028.1381, 1028.0851, 1028.0331, 1027.9827, 1027.9285, 1027.8749, 1027.8214, 1027.7714, 1027.7135, 1027.653, 1027.5984, 1027.5464, 1027.4911, 1027.4349, 1027.3798, 1027.3098, 1027.2406, 1027.1884, 1027.1222, 1027.0693, 1027.0184, 1026.9578, 1026.9069, 1026.8369, 1026.7656, 1026.6857, 1026.5956, 1026.4814, 1026.3639, 1026.263, 1026.0757, 1025.9543, 1025.7444, 1025.5826, 1025.4564, 1025.359, 1025.2089, 1025.1049, 1024.9454, 1024.7924, 1024.6616, 1024.5201, 1024.4451, 1024.2979, 1024.1198, 1024.0754, 1024.0515, 1024.032, 1024.0106, 1023.986, NaN, NaN, 1029.2056, 1029.1726, 1029.1321, 1029.0793, 1029.0192, 1028.9631, 1028.9062, 1028.8542, 1028.8013, 1028.7496, 1028.6981, 1028.6461, 1028.595, 1028.5399, 1028.4784, 1028.4246, 1028.3636, 1028.3114, 1028.257, 1028.1968, 1028.149, 1028.095, 1028.0413, 1027.9828, 1027.9247, 1027.8691, 1027.8184, 1027.7631, 1027.7002, 1027.6339, 1027.5648, 1027.4984, 1027.4387, 1027.3729, 1027.301, 1027.229, 1027.1539, 1027.0767, 1027.001, 1026.9393, 1026.8689, 1026.7963, 1026.7273, 1026.6482, 1026.5535, 1026.4492, 1026.3112, 1026.1482, 1025.9958, 1025.87, 1025.7032, 1025.6229, 1025.5226, 1025.4124, 1025.309, 1025.2014, 1025.1244, 1025.0151, 1024.831, 1024.7183, 1024.6432, 1024.5609, 1024.4564, 1024.2938, 1024.1024, 1024.0723, 1024.0459, 1024.0248, 1024.0123, NaN, NaN, 1029.1824, 1029.1532, 1029.1149, 1029.069, 1029.0289, 1028.9807, 1028.935, 1028.887, 1028.8392, 1028.7882, 1028.7339, 1028.6891, 1028.6416, 1028.5895, 1028.5372, 1028.4893, 1028.4387, 1028.3883, 1028.3401, 1028.2903, 1028.2407, 1028.1891, 1028.1372, 1028.0862, 1028.027, 1027.9719, 1027.918, 1027.8624, 1027.8201, 1027.7698, 1027.7218, 1027.6722, 1027.6183, 1027.5647, 1027.5042, 1027.4469, 1027.3888, 1027.3246, 1027.2627, 1027.1951, 1027.1185, 1027.0518, 1026.9684, 1026.8843, 1026.8002, 1026.7164, 1026.6168, 1026.5316, 1026.3953, 1026.2765, 1026.1641, 1026.0345, 1025.8661, 1025.6985, 1025.5651, 1025.4205, 1025.3138, 1025.2013, 1025.0809, 1024.9442, 1024.8096, 1024.6882, 1024.5729, 1024.4539, 1024.183, 1024.1042, 1024.0608, 1024.0361, 1024.0112, 1023.33923, 1022.77374, 1022.87177, NaN, NaN, 1027.1027, 1027.0527, 1026.9895, 1026.8816, 1026.8083, 1026.7448, 1026.6655, 1026.5532, 1026.4542, 1026.4225, 1026.3198, 1026.0619, 1026.3538, 1026.2589, 1026.2379, 1026.1927, 1026.0197, 1026.5497, 1028.2483, 1028.1919, 1028.1349, 1028.0778, 1028.0194, 1027.9597, 1027.895, 1027.8373, 1027.79, 1027.7281, 1027.6746, 1027.6151, 1027.5662, 1027.5098, 1027.4513, 1027.3838, 1027.325, 1027.2604, 1027.1897, 1027.111, 1027.0371, 1026.9642, 1026.8978, 1026.8147, 1026.7201, 1026.6237, 1026.4954, 1026.287, 1026.1293, 1026.0052, 1025.8566, 1025.7249, 1025.5902, 1025.4452, 1025.3221, 1025.1984, 1025.083, 1024.9622, 1024.7975, 1024.6351, 1024.537, 1024.2335, 1024.1045, 1024.0698, 1024.0321, 1023.99316, 1023.918, 1023.87006, 1023.85315, NaN, NaN, 1029.1819, 1029.1543, 1029.1207, 1029.0773, 1029.0374, 1028.9895, 1028.938, 1028.8892, 1028.8445, 1028.7977, 1028.7533, 1028.7012, 1028.6469, 1028.5953, 1028.5454, 1028.4901, 1028.4358, 1028.3768, 1028.3225, 1028.2682, 1028.2158, 1028.1595, 1028.102, 1028.0414, 1027.9855, 1027.9337, 1027.8846, 1027.8323, 1027.774, 1027.7223, 1027.6632, 1027.6145, 1027.5653, 1027.5105, 1027.4536, 1027.3982, 1027.3367, 1027.2698, 1027.2148, 1027.1434, 1027.0583, 1026.9688, 1026.8986, 1026.8114, 1026.7194, 1026.6346, 1026.5344, 1026.4172, 1026.2883, 1026.1625, 1026.0048, 1025.8265, 1025.6823, 1025.5494, 1025.4243, 1025.2777, 1025.1685, 1025.0848, 1024.9729, 1024.8093, 1024.6874, 1024.5876, 1024.4196, 1024.1211, 1024.0579, 1024.0299, 1023.9956, 1023.9496, 1023.8636, 1023.8369, NaN, NaN, 1029.2056, 1029.1698, 1029.1311, 1029.0841, 1029.034, 1028.9757, 1028.9218, 1028.8751, 1028.8229, 1028.765, 1028.7142, 1028.6672, 1028.6173, 1028.5658, 1028.5121, 1028.4548, 1028.3873, 1028.3318, 1028.2836, 1028.2334, 1028.186, 1028.1364, 1028.0844, 1028.0265, 1027.9681, 1027.9054, 1027.8444, 1027.7909, 1027.7362, 1027.6774, 1027.616, 1027.5663, 1027.5187, 1027.4633, 1027.3944, 1027.3296, 1027.2681, 1027.2109, 1027.151, 1027.0874, 1027.0145, 1026.9387, 1026.8582, 1026.7465, 1026.6467, 1026.5366, 1026.3909, 1026.2695, 1026.1509, 1026.0287, 1025.8768, 1025.6686, 1025.4951, 1025.3572, 1025.255, 1025.1534, 1025.062, 1024.9601, 1024.8486, 1024.718, 1024.561, 1024.3793, 1024.1031, 1024.0652, 1024.0062, 1023.9654, 1023.87146, 1023.76965, 1023.7216, 1023.7038, NaN, NaN, 1029.1951, 1029.1686, 1029.1338, 1029.084, 1029.0255, 1028.9711, 1028.9149, 1028.8619, 1028.8079, 1028.7574, 1028.706, 1028.6536, 1028.6033, 1028.5447, 1028.4911, 1028.4344, 1028.384, 1028.3314, 1028.2836, 1028.2255, 1028.1709, 1028.1116, 1028.0555, 1027.9834, 1027.9183, 1027.859, 1027.8048, 1027.7446, 1027.6831, 1027.6194, 1027.5607, 1027.5001, 1027.45, 1027.3882, 1027.3225, 1027.2614, 1027.1863, 1027.1002, 1027.0404, 1026.9794, 1026.9146, 1026.8278, 1026.7101, 1026.5908, 1026.4713, 1026.3269, 1026.1584, 1026.0688, 1025.8171, 1025.6188, 1025.4681, 1025.3152, 1025.1962, 1025.0707, 1024.9707, 1024.8568, 1024.716, 1024.5524, 1024.2819, 1024.0677, 1024.0024, 1023.91315, 1023.85223, 1023.7871, 1023.7425, 1023.70294, 1023.6669, NaN, NaN, 1029.2183, 1029.1901, 1029.1539, 1029.1084, 1029.0638, 1029.0116, 1028.9596, 1028.9114, 1028.858, 1028.8073, 1028.7563, 1028.7057, 1028.6564, 1028.6085, 1028.5544, 1028.5062, 1028.4521, 1028.3926, 1028.3458, 1028.2966, 1028.2467, 1028.199, 1028.1526, 1028.1052, 1028.0509, 1027.9956, 1027.9368, 1027.8784, 1027.8243, 1027.7795, 1027.7284, 1027.6572, 1027.5887, 1027.5345, 1027.4811, 1027.4288, 1027.3741, 1027.3235, 1027.2705, 1027.2048, 1027.134, 1027.0597, 1026.9883, 1026.9156, 1026.8177, 1026.7164, 1026.632, 1026.5442, 1026.4297, 1026.3182, 1026.2056, 1026.0596, 1025.9408, 1025.6888, 1025.5078, 1025.3514, 1025.2622, 1025.1376, 1025.0498, 1024.948, 1024.794, 1024.5989, 1024.3362, 1024.0897, 1024.0116, 1023.9668, 1023.94556, 1023.90814, 1023.8532, 1023.7462, 1023.69745, NaN, NaN, 1029.1979, 1029.1714, 1029.1365, 1029.0914, 1029.0492, 1029.0062, 1028.9557, 1028.9132, 1028.8625, 1028.809, 1028.7599, 1028.7117, 1028.6705, 1028.627, 1028.5742, 1028.5288, 1028.4797, 1028.4315, 1028.3851, 1028.3367, 1028.2853, 1028.2397, 1028.1946, 1028.1538, 1028.1062, 1028.0554, 1027.9978, 1027.9537, 1027.8994, 1027.8463, 1027.7933, 1027.7396, 1027.6923, 1027.6405, 1027.583, 1027.5208, 1027.469, 1027.4146, 1027.353, 1027.2911, 1027.2324, 1027.1733, 1027.113, 1027.0535, 1026.9913, 1026.929, 1026.8536, 1026.7533, 1026.6653, 1026.5682, 1026.4741, 1026.3558, 1026.2263, 1026.1129, 1026.0022, 1025.9304, 1025.8315, 1025.6974, 1025.5515, 1025.4197, 1025.3068, 1025.1886, 1025.0574, 1024.9268, 1024.8187, 1024.6147, 1024.3414, 1024.0525, 1023.9776, 1023.9523, 1023.92487, 1023.89343, 1023.8251, NaN, NaN, 1029.2056, 1029.1742, 1029.1393, 1029.0859, 1029.0317, 1028.9747, 1028.9204, 1028.8667, 1028.8103, 1028.7559, 1028.6996, 1028.6473, 1028.593, 1028.5374, 1028.4802, 1028.4243, 1028.37, 1028.318, 1028.266, 1028.2146, 1028.1649, 1028.1084, 1028.0559, 1028.0072, 1027.9619, 1027.9113, 1027.8599, 1027.7998, 1027.7404, 1027.688, 1027.6437, 1027.5951, 1027.5249, 1027.4681, 1027.4132, 1027.3536, 1027.3026, 1027.2546, 1027.1908, 1027.1161, 1027.0364, 1026.9498, 1026.867, 1026.772, 1026.6616, 1026.5334, 1026.4338, 1026.3196, 1026.2236, 1026.1035, 1025.9862, 1025.8441, 1025.7045, 1025.5632, 1025.4058, 1025.3165, 1025.201, 1025.0951, 1024.9543, 1024.8737, 1024.7563, 1024.5712, 1024.3878, 1024.065, 1024.0044, 1023.9719, 1023.94025, 1023.90027, 1023.8211, 1023.7925, NaN, NaN, 1029.2107, 1029.1825, 1029.1456, 1029.0908, 1029.0342, 1028.9812, 1028.9293, 1028.8787, 1028.8252, 1028.7767, 1028.7279, 1028.6759, 1028.6249, 1028.5767, 1028.5239, 1028.4719, 1028.4236, 1028.3696, 1028.3108, 1028.2592, 1028.1973, 1028.1422, 1028.089, 1028.0295, 1027.975, 1027.9126, 1027.8505, 1027.7845, 1027.7087, 1027.6478, 1027.5828, 1027.5062, 1027.4321, 1027.3774, 1027.3102, 1027.2441, 1027.1736, 1027.1053, 1027.0331, 1026.9603, 1026.8815, 1026.8087, 1026.696, 1026.5579, 1026.4458, 1026.2793, 1026.1268, 1025.9608, 1025.8234, 1025.6335, 1025.4741, 1025.3484, 1025.255, 1025.1116, 1024.9703, 1024.8705, 1024.78, 1024.5677, 1024.428, 1024.3308, 1024.1941, 1024.1184, 1024.0305, 1023.92395, 1023.8574, 1023.8284, 1023.81354, NaN, NaN, 1029.2263, 1029.1989, 1029.1608, 1029.1104, 1029.0594, 1029.0042, 1028.9478, 1028.8899, 1028.8392, 1028.7836, 1028.7269, 1028.6747, 1028.6241, 1028.5739, 1028.517, 1028.4675, 1028.4161, 1028.365, 1028.3143, 1028.2607, 1028.2036, 1028.1466, 1028.0956, 1028.0438, 1027.9943, 1027.9419, 1027.8855, 1027.8328, 1027.7831, 1027.7205, 1027.6604, 1027.6118, 1027.5619, 1027.5023, 1027.4459, 1027.3777, 1027.3171, 1027.2496, 1027.1898, 1027.1165, 1027.0404, 1026.9624, 1026.8827, 1026.786, 1026.6906, 1026.5563, 1026.3823, 1026.1809, 1026.0239, 1025.8798, 1025.7681, 1025.6389, 1025.5059, 1025.3774, 1025.2712, 1025.156, 1025.0128, 1024.9073, 1024.7926, 1024.6017, 1024.4636, 1024.3448, 1024.2166, 1024.0723, 1024.0038, 1023.96277, 1023.91876, 1023.8949, NaN, NaN, 1029.2084, 1029.178, 1029.1422, 1029.09, 1029.0332, 1028.9755, 1028.9247, 1028.8672, 1028.8098, 1028.7567, 1028.7013, 1028.6454, 1028.5933, 1028.544, 1028.4922, 1028.4386, 1028.3895, 1028.3383, 1028.2869, 1028.2349, 1028.1881, 1028.139, 1028.0853, 1028.0333, 1027.9761, 1027.9083, 1027.8602, 1027.8088, 1027.7542, 1027.6927, 1027.6393, 1027.581, 1027.5237, 1027.4652, 1027.402, 1027.3381, 1027.2797, 1027.1953, 1027.1194, 1027.0626, 1026.9966, 1026.921, 1026.8406, 1026.752, 1026.6407, 1026.5421, 1026.3978, 1026.2273, 1026.0791, 1025.928, 1025.7864, 1025.6555, 1025.564, 1025.4584, 1025.3256, 1025.2289, 1025.141, 1025.0697, 1024.9724, 1024.8483, 1024.683, 1024.6154, 1024.4935, 1024.31, 1024.1628, 1024.0841, 1023.9737, 1023.92755, 1023.8968, NaN, NaN, 1029.2197, 1029.1919, 1029.1571, 1029.1085, 1029.0615, 1029.0137, 1028.9609, 1028.9119, 1028.8615, 1028.8104, 1028.7607, 1028.712, 1028.6602, 1028.6062, 1028.5527, 1028.4995, 1028.4475, 1028.3938, 1028.3397, 1028.2899, 1028.2401, 1028.1837, 1028.1327, 1028.0789, 1028.0189, 1027.9559, 1027.9095, 1027.8551, 1027.8005, 1027.7511, 1027.6978, 1027.6477, 1027.5968, 1027.5488, 1027.508, 1027.4517, 1027.4075, 1027.3417, 1027.2758, 1027.2189, 1027.1566, 1027.0859, 1027.038, 1026.9708, 1026.9147, 1026.8014, 1026.6995, 1026.5732, 1026.4589, 1026.3197, 1026.1748, 1026.0334, 1025.9116, 1025.779, 1025.6469, 1025.5505, 1025.4602, 1025.3309, 1025.235, 1025.1748, 1025.0845, 1024.9647, 1024.8716, 1024.7539, 1024.6245, 1024.5116, 1024.3785, 1024.1409, 1023.9984, 1023.9596, 1023.9343, 1023.91833, NaN, NaN, 1029.2227, 1029.1931, 1029.152, 1029.1008, 1029.0542, 1029.0039, 1028.9434, 1028.8835, 1028.8262, 1028.7737, 1028.7195, 1028.6617, 1028.6053, 1028.5463, 1028.4886, 1028.428, 1028.3755, 1028.3228, 1028.2747, 1028.2197, 1028.1692, 1028.1193, 1028.0651, 1028.0183, 1027.9626, 1027.9158, 1027.8651, 1027.8063, 1027.7502, 1027.6962, 1027.6409, 1027.5836, 1027.5298, 1027.467, 1027.3909, 1027.3342, 1027.2731, 1027.2091, 1027.146, 1027.0762, 1027.0048, 1026.9347, 1026.833, 1026.7405, 1026.6241, 1026.5162, 1026.3948, 1026.2491, 1026.1381, 1025.9296, 1025.7224, 1025.6196, 1025.4938, 1025.4197, 1025.3538, 1025.2363, 1025.1388, 1025.0667, 1024.9775, 1024.8593, 1024.7313, 1024.5498, 1024.4442, 1024.2716, 1024.0798, 1024.0043, 1023.96027, 1023.9362, 1023.911, 1023.8951, NaN, NaN, 1029.2385, 1029.2089, 1029.1733, 1029.1277, 1029.0776, 1029.028, 1028.9784, 1028.93, 1028.8794, 1028.8315, 1028.7839, 1028.7307, 1028.6754, 1028.6248, 1028.5715, 1028.5227, 1028.4698, 1028.4155, 1028.3661, 1028.3159, 1028.2601, 1028.2039, 1028.1484, 1028.0868, 1028.0288, 1027.9717, 1027.909, 1027.8524, 1027.8, 1027.7494, 1027.6897, 1027.637, 1027.5771, 1027.5186, 1027.4675, 1027.4135, 1027.353, 1027.2964, 1027.2413, 1027.1829, 1027.1149, 1027.0338, 1026.9543, 1026.8577, 1026.766, 1026.6893, 1026.5865, 1026.4818, 1026.3145, 1026.1715, 1026.0026, 1025.8903, 1025.7388, 1025.5305, 1025.3928, 1025.2631, 1025.1276, 1025.04, 1024.9138, 1024.7927, 1024.6299, 1024.4224, 1024.218, 1024.0759, 1024.0306, 1024.0013, 1023.9687, 1023.92957, 1023.8957, 1023.8821, NaN, NaN, 1029.2394, 1029.2128, 1029.1753, 1029.1293, 1029.0798, 1029.0306, 1028.9728, 1028.9232, 1028.8695, 1028.817, 1028.7623, 1028.7019, 1028.6409, 1028.582, 1028.5295, 1028.4779, 1028.426, 1028.369, 1028.3099, 1028.2556, 1028.2025, 1028.145, 1028.0924, 1028.0372, 1027.9794, 1027.9216, 1027.8645, 1027.8064, 1027.7513, 1027.6945, 1027.6312, 1027.5757, 1027.5223, 1027.4672, 1027.4062, 1027.3353, 1027.271, 1027.1997, 1027.1212, 1027.0383, 1026.9407, 1026.8539, 1026.7537, 1026.6069, 1026.4542, 1026.2913, 1026.1257, 1026.0177, 1025.937, 1025.8104, 1025.6943, 1025.5299, 1025.4039, 1025.2909, 1025.1569, 1025.058, 1024.9913, 1024.8665, 1024.6887, 1024.436, 1024.2517, 1024.111, 1024.0791, 1024.0537, 1024.0128, 1023.93823, 1023.88947, 1023.8679, NaN}
    DOXY = 
      {NaN, 31.683392429188327, 31.347443551015285, 31.969393597180186, 32.69823186866394, 33.39011221503253, 33.97048544798978, 34.66100612930025, 35.42510375960818, 36.152835963468824, 37.175658636808016, 38.3090202457831, 39.516021954528505, 41.130667137281684, 43.111816837953064, 44.83326897290415, 46.59196455395993, 49.051064811438955, 51.76656043421727, 54.00058745598457, 56.45904409434231, 58.62482057435487, 59.5079467031923, 59.28790113637347, 60.61049734714558, 64.42199412341932, 65.2319680517248, 67.42497517157713, 67.86400601068829, 68.01416983772687, 71.54368073885168, 74.34324356496539, 72.28630417430776, 72.35167752538827, 73.8221462951993, 74.25747563477601, 76.01913082864766, 78.8836872689865, 84.24609203359223, 82.99563339671371, 83.4273967415388, 85.253460173305, 85.97387993274484, 87.61476872412081, 90.3712316913608, 92.76772277445262, 94.78746319763066, 98.27637857627079, 105.81487608002497, 115.57447517700233, 129.41550172121242, 142.32134510801689, 154.71284205502243, 173.6099672443893, 190.8576908893167, 204.29160937096665, 215.33521705719852, 224.77129403627757, 233.3820555964706, 242.48310414816578, 250.51432381651438, 257.54355266561925, 264.88540864468183, 274.5623378245004, 275.0770201129301, 257.6481454624237, 250.02699812373055, 249.6864036141998, 250.0931833767521, 250.0694516971574, 249.49344194481665, 249.10359267546377, NaN, NaN, 31.31497106272985, 30.941832175764592, 31.52721961552659, 32.1815113540639, 32.946509867851795, 33.63536206505905, 34.25062720199403, 35.086644273305154, 36.292229534487184, 37.79190840349752, 39.550585235273424, 41.232939257016184, 42.87816698240942, 44.81861814131099, 46.6465043310144, 48.47539540362197, 50.04294079562156, 51.9073026407083, 54.509983756708074, 57.69935857808647, 60.66893610757869, 62.93611763753828, 64.18027106365297, 64.2481901171757, 65.27817492231465, 67.48231534859926, 69.6856636875284, 69.45536327847782, 65.34616918604912, 67.11981304022575, 74.54069651825499, 76.74464815522965, 74.76525686730064, 74.17747357091697, 76.74074431153977, 78.06395162109665, 78.50630318219102, 80.85875600269694, 82.31928386318548, 83.4816493822829, 85.97143032773602, 87.43080304623334, 89.6233727019703, 92.56488813798097, 95.14178473516841, 99.1950518425506, 104.88689808169852, 112.98875018667114, 126.44133035358199, 149.00119590701138, 170.23318817442092, 190.10800629860265, 210.30954677743995, 222.92844671703622, 233.73858437439415, 238.8215942456326, 243.8921807484052, 255.33621788386995, 261.2093836690566, 265.8024614796466, 262.54134889001506, 248.58201127237754, 247.35170405815705, 248.06511793525982, 247.88260893068338, 247.17303933536087, 247.15290491358218, NaN, NaN, 30.31556174087382, 29.722518532564855, 30.56756564318249, 31.4446973098675, 32.58233275004621, 33.60627921577216, 34.55595258842796, 35.32039071661771, 36.49138668351489, 37.69891027188058, 39.49641446784758, 41.58944711352048, 43.7911312437416, 45.40130986184979, 46.97377479416805, 48.655966835671045, 50.411654391808426, 52.27540223863598, 54.88275790194432, 57.59423053071894, 58.753613495294225, 59.61928469612495, 61.37310136816033, 64.74890014675964, 68.0450483203491, 70.23473373810599, 73.7598471967512, 75.96841763463632, 76.99172878665878, 77.364538655341, 73.03751708033275, 69.59075388872056, 70.10707648642331, 72.31746787367626, 73.93527429358387, 74.00465407286954, 76.58068565695396, 81.51511949544762, 84.0876383015575, 85.18748107936595, 87.26997721601346, 89.28011858375955, 89.827321634716, 92.21677776990505, 92.3999024171428, 94.05522891155617, 102.34045370152903, 109.67814384541234, 112.96256116291742, 114.77547177083878, 122.71995508834924, 140.44490035910422, 150.39121925665697, 169.47257517913562, 183.11015507992363, 198.03952171220888, 211.87394146367498, 224.3143290764998, 234.69665480684063, 240.02331961581527, 244.17013117891744, 256.81341039785286, 263.78866844276047, 251.04708248531946, 248.23730414535297, 247.2554471453139, 245.8263518579726, 245.800822047414, 246.03869315288145, 246.29884987595224, NaN, NaN, 32.910008922834784, 32.27833568680218, 32.90027110242337, 34.44370899284209, 35.43011283270054, 36.60132057553497, 37.585508525715156, 39.19979632584583, 40.663932608495756, 43.16475010594799, 45.77248144368395, 47.971963394456296, 49.98531332429777, 51.777174930150636, 53.34626670863937, 55.21096577445153, 57.18536719369933, 59.603171643764476, 61.4260686957624, 62.25272360542857, 63.71152530382979, 65.97555849903092, 67.35437354740706, 69.02981408006956, 71.29174861118999, 75.10421077448133, 80.46225071964868, 83.99429695181863, 80.40127171626308, 77.24113824557304, 75.8701350518854, 73.68591705281598, 75.30820347651454, 76.2654146629525, 77.58961620011442, 79.93146638409364, 82.19637358122317, 83.28549437918714, 84.67703958955084, 87.2406196232687, 87.95771124422374, 88.49461964637531, 89.76766258928969, 91.59162353713414, 93.78340852345349, 97.6361691898264, 104.98450976201619, 113.44725257449743, 128.9317446944312, 142.948236148521, 157.1774268410845, 178.6666286028305, 198.37176797283797, 218.1026313980898, 234.53625692765286, 243.63788194642797, 247.12171852770877, 253.34308061892833, 265.02566366783924, 264.21654944877986, 246.7916976060655, 243.9165772364817, 244.17990140092138, 244.57699700213743, 244.83688699886721, NaN, NaN, 31.388444606774023, 30.64604864783854, 31.046329408026544, 32.44257928697277, 34.318007651751024, 36.154249411799746, 37.767521663041144, 39.41833302490893, 41.401539692105224, 43.198394015520975, 45.55070276007592, 47.715683663165684, 49.95386163030589, 52.117783790807, 53.35548454570277, 54.33485992889705, 55.46202880417194, 56.47850427134795, 58.86549920752095, 60.69050940469694, 62.29687242263562, 63.973614374498766, 65.57498982474965, 66.66139679672379, 68.55737120094737, 70.22867390134104, 72.12148302674878, 75.63791599752734, 81.88691477758167, 84.77027235107663, 80.54433414358333, 78.15905239835796, 77.20872981249245, 75.59300066076466, 76.76481885637973, 78.22182880554364, 79.45965087553884, 80.9921574557938, 82.52182289274901, 83.38767803109407, 84.47456567842417, 85.12245182523141, 86.43752157871091, 87.30988263517229, 88.62371187151605, 90.81419068475779, 93.00503639466717, 96.30125758082741, 102.71035592521787, 109.54923749615021, 121.92634232198147, 138.5229999164271, 157.16785029460158, 181.6413988250454, 199.9146080498324, 210.42466661463533, 223.80297840625494, 237.73110035252586, 247.79748478236974, 263.39872852026207, 267.63376232555214, 250.58958734893764, 244.89371022182192, 245.00782144520352, 244.95130147231802, 245.1162269634463, 245.3664201207841, 245.629311073959, NaN, NaN, 31.165726826835012, 30.127472447862615, 30.639046312061673, 31.36794907332996, 32.3937467725737, 33.6777166867089, 35.47867193128366, 37.20382933152928, 38.81845398617741, 41.245825298405606, 43.63468573468178, 45.837789147417396, 48.26331119790948, 49.83487257065503, 51.85220587632646, 53.49934842692196, 55.476707398349824, 56.456724714551825, 57.399800856136785, 59.41771773396418, 61.72525083642554, 63.108452067793024, 65.37666046808954, 66.092169645594, 68.51171950187965, 72.0304497190015, 74.66140369556703, 77.58820335885785, 82.36600812358118, 83.36610138148262, 77.39748597660378, 75.41998933221203, 75.27504267345444, 74.67543202270976, 75.03369411837859, 76.49424949619487, 78.63030867638564, 80.90472257352845, 82.51268181981351, 83.38095104624018, 84.28389187074151, 85.29835016360396, 85.7964647845166, 86.56304648394739, 85.77941321072458, 88.8529935054288, 89.09900573213515, 88.57321839680867, 90.10009041278784, 93.68660627893696, 98.81681352594542, 101.89916148893134, 104.45642097701483, 106.50295212751085, 115.79657495910524, 139.82542723131175, 170.4387365595193, 193.83045049211714, 212.98414646768427, 230.09821507418664, 241.05917582350034, 250.54444162180582, 262.83510071747804, 270.6890514906187, 270.9568433384986, 257.91676053576333, 247.93524021330137, 246.46349804791296, 244.27575075215842, 243.91501708244596, 244.0884415393821, 244.2730740840563, NaN, NaN, 31.055557630507835, 30.202456385934504, 30.714434627612746, 31.814673304653496, 33.32041067879863, 35.232593343898145, 36.844989628312554, 37.60786159985361, 39.22140125162537, 40.3892211763562, 41.92858751664428, 45.205075189899745, 48.217679605565536, 50.52909928381305, 52.54221141676462, 54.002597973671925, 55.5357760069679, 57.14289152187621, 58.861726248962064, 61.280480654254504, 62.43998218620632, 64.48781335442095, 66.23606270257339, 68.72523474772474, 70.98608181922854, 72.06866460468618, 74.92534596823758, 79.61817268826105, 82.8503836327882, 84.17579615582795, 81.3470998834181, 75.38640744393778, 74.88380565673353, 75.1044992782121, 75.980278863568, 77.21794773740885, 79.50903084225178, 82.0025543933607, 83.31612816711687, 84.40268474829308, 85.01103520947233, 85.87420591052633, 86.15893762352674, 85.26513094830894, 86.71859434984948, 87.8768522135614, 89.32632029604173, 89.3119563430859, 91.06134851029923, 98.68289251515185, 102.19071455420162, 104.82362084382383, 109.82836448818728, 127.83942034600415, 163.96088911412744, 193.08074375963375, 214.62418089579535, 232.14279440614604, 239.95378518389865, 248.56798010542718, 260.1810175465726, 267.38753581497315, 261.8861878167376, 249.39311979198945, 244.58422135796278, 243.46451528846126, 243.75340449767086, 244.041420280437, 244.23210814712255, NaN, NaN, 33.64594586289366, 32.24044577760941, 32.899344942269934, 34.14746136666166, 35.802947823914124, 37.157933689795065, 38.62549320035493, 40.31363598242659, 42.07498386794718, 43.02008585238358, 44.671499138852944, 46.763793885342636, 48.89125381871034, 51.316986683000906, 53.627062486837175, 55.30935540405026, 56.80605027145806, 58.48767454466596, 60.093887798973874, 61.32817946500989, 62.491327510514495, 65.72082193784136, 67.02367145931584, 68.32937325907345, 70.30025481122219, 73.08191725706718, 78.07583233195511, 81.82642498112675, 80.81287035596736, 80.16082259355316, 77.76321738058729, 75.12585089100098, 74.68255751771396, 75.34180415480185, 76.14539822544161, 76.58051869632857, 77.98533792530888, 79.67635499435191, 80.6189314280156, 82.07674950511115, 83.27596218271424, 84.43843641217671, 85.30753785572746, 85.59030056346128, 85.58028725312109, 85.85637242321437, 89.07080957543725, 88.7592135102645, 89.33104602599846, 92.55116635332568, 97.83597462299271, 102.23121300183179, 103.97358107191478, 106.01869878381336, 113.67749285033987, 140.57570114849455, 174.93337357949184, 196.0145911066971, 215.18661803212268, 231.8575963715913, 244.31815687570491, 255.5055769689811, 262.4369324140268, 265.82204942086054, 248.45508096927892, 243.0642997304313, 243.5777700139025, 244.0879678442, 244.43537491770888, NaN, NaN, 45.15980647727301, 34.080872460515955, 33.0787629889868, 33.844594685675865, 35.38620102571013, 36.260713208373495, 37.134228192532234, 38.121082380121926, 40.328114782814716, 42.97648701096595, 45.068803162851545, 46.494965584002685, 48.144196267853395, 50.34621745472326, 51.99183626274744, 54.08345309228603, 56.06139518208326, 57.927904720792235, 59.90403897565767, 61.437303312861424, 62.748317071870055, 65.05558127690125, 67.13674465006093, 69.29285644938312, 72.11097686101967, 75.18792987296752, 79.73675105727237, 82.68521791402335, 81.77281410713148, 78.4394057190174, 77.31386087864668, 76.43722065256722, 75.66824789310398, 75.82440604744359, 76.0413487122382, 77.55217126075397, 79.90050103843059, 81.28987166304927, 82.89808012120282, 84.13178923847832, 85.14337406658527, 85.79409806260752, 86.6585039019304, 87.96232056911062, 88.60807505093618, 88.59072516845339, 89.90434949230372, 91.88054669775947, 94.07692290853046, 97.38282439500998, 104.01138466486113, 110.18730445232579, 117.03020105480103, 131.41642941721753, 155.39890966086875, 180.57636161543803, 200.69312637770355, 220.32393918610214, 231.82880330533874, 240.7786583691914, 247.23979583534796, 256.07979878678105, 259.4982707401744, 267.5696239944786, 272.29591771214893, 265.50444918451547, 252.4400833625959, 247.15492259855642, 245.04346709562836, 244.92175466282558, 244.9971006350824, 245.18530339886354, NaN, NaN, 34.823029933665545, 31.64402807335673, 31.785431259694423, 32.848229103571704, 34.0949846586896, 35.37597206047416, 36.54587498901889, 37.78938153248042, 39.03200051574412, 40.20149345335639, 41.888220514124, 43.905891186763625, 45.73683466793086, 47.34580310592165, 48.77020359976682, 50.71323811072122, 53.022825280619195, 55.777408823157735, 58.67573505060181, 60.50084909936472, 62.84398565252563, 65.07172875912887, 66.67174309571917, 69.41531221217024, 73.1168334440458, 76.48395161803285, 79.64027225727115, 80.85403795162372, 78.3056190345604, 75.2250149840704, 74.23646898796136, 73.02647317009026, 76.0041958222451, 77.37235545079834, 77.46994814458596, 78.15720033534384, 81.01896310120361, 83.25285522527463, 84.23047107662386, 85.0558106840188, 85.8471160496729, 86.49491111753775, 88.25069327127656, 89.78387697036328, 91.98072498488943, 97.05335606284655, 103.22233179564049, 109.61711638356658, 121.5487797194495, 136.3889034216868, 161.92046531463353, 180.38556975526643, 204.13664560343665, 222.56093944542968, 231.6075732874091, 240.48039784158868, 247.0749171861981, 252.52642671719434, 260.17707770995617, 267.52549768980947, 266.5741233930188, 256.81618011913474, 252.75992300987926, 249.01370047440903, 248.45607600660702, 248.6488560275085, NaN, NaN, 51.91673017421926, 35.67121821244097, 33.74526499746066, 34.03153784474652, 34.75976482719067, 35.78434063178029, 37.40008212143278, 38.717094793935495, 40.03604175151854, 41.944593897944465, 43.55521174683102, 45.16849325218967, 47.223498756793134, 49.12766854070001, 51.0294319652065, 52.193721196478656, 53.95030716362958, 56.88962116973497, 59.37844235486433, 60.9825153605851, 63.73195615986454, 65.73625873986622, 67.93020150831974, 70.6716000511623, 74.09075116337861, 76.06990997166824, 77.69329046800765, 77.5466936850165, 73.91649173152746, 72.23191703412787, 72.7156572623685, 72.11999962315295, 73.21671586751698, 76.30560724581954, 77.43744492201851, 77.95227306845146, 79.15649275704854, 81.49883366812499, 82.3718930266646, 84.97169631803337, 86.39141463741687, 87.84942292211029, 90.04005428188965, 90.94209843575608, 91.48953214062183, 90.9322405104939, 94.97126180466384, 99.73992254302767, 106.1739054929728, 117.757228541104, 131.04445202812033, 146.7510013140898, 167.4589515334269, 184.54586923366142, 204.51683608509472, 218.54176569951528, 227.15748640787217, 236.12319271471645, 245.79807978568712, 251.32985456325977, 258.8218101676789, 266.86751099842974, 267.3241683588136, 263.63913985980633, 257.5592947661353, 252.08619066964883, 250.98568746472344, 251.09157766731855, NaN, NaN, 32.50329625064442, 32.24033204794143, 32.82527551995867, 33.59117110763454, 34.43105527659845, 35.45465203236205, 36.58802743563318, 37.68482070651241, 39.00123901778322, 40.133649090762894, 41.56071163804159, 43.02414227695593, 44.524326080032765, 46.17121034563424, 48.00279373850686, 49.86948263556187, 51.88462785084255, 54.59896327080189, 57.34925224840809, 60.46861464022525, 63.290813907061256, 66.07547925705535, 68.67324897569618, 70.79496241046401, 72.0751577663838, 72.36789285033153, 75.49510585769536, 75.5424102889436, 71.32955607000488, 73.75566944515388, 73.69700073181657, 74.65389413701503, 76.52194538925083, 77.4798572246344, 78.43775788981429, 80.74678235273211, 81.69498712513261, 83.0840886927445, 85.27493957981012, 85.92100067341111, 86.71456518728449, 87.98782388640367, 87.61170451226963, 88.33756743712411, 88.14446978168583, 89.05345905167843, 94.74126315935219, 102.45334394344204, 108.14789490534874, 116.61821868212941, 130.0944831120008, 147.08884429637018, 167.80125725265574, 185.44531150605118, 208.64306259790442, 222.6742767897797, 229.04074068163806, 236.2693706495072, 244.25513054605588, 250.33863979065515, 255.44911420509186, 260.7929109601348, 264.0509445608782, 261.5444479832838, 257.7377013516262, 254.7031266934265, 251.21491957859638, 250.60914143285422, 251.01442761408413, NaN, NaN, 36.01215428696288, 33.53452485923902, 33.601529449940706, 34.405038421670824, 34.87560965154473, 35.78944456779221, 36.591244936157516, 37.46698536880114, 38.2687760058943, 39.40188776594399, 40.57133286126466, 41.92589734956759, 43.427255262804934, 44.92751356066545, 46.35320925844171, 48.29600118802958, 50.5325828683771, 52.73085784565606, 55.33422058528008, 57.899413705068156, 60.836055718829854, 64.02848539623629, 66.85013955452219, 69.08522716313261, 69.88432970420531, 71.57454148131919, 72.45445175081491, 73.15112147479427, 72.42164103087808, 70.70794520802306, 71.70817495727586, 72.437354704102, 72.20995150093607, 72.76131167471725, 74.5271503163428, 76.58587635592468, 76.84601033520516, 78.15790721640485, 79.43472873973072, 80.56895950799893, 81.58900650949039, 83.78580640854834, 86.3462537132745, 86.33275553241828, 86.68341147502379, 86.85032099485177, 88.12728552423565, 90.69632319852126, 94.17975875043875, 98.76953401648942, 105.75394793587024, 113.67237939345036, 125.09512958893275, 145.79471696414524, 166.28403143805988, 179.96495445399614, 197.68974775306162, 216.80314391434817, 229.57675776162927, 240.07641963943018, 248.964840118762, 256.74411959699796, 262.0687165021344, 268.21047086443417, 265.672171377732, 258.591468692651, 252.65840281017708, 250.5005005561584, 250.17975657408272, NaN, NaN, 38.52425767007105, 34.754071046445155, 34.78434386587644, 35.587439245432854, 36.86817861869674, 37.741223856965604, 38.31801991369174, 39.56175971628323, 40.98867507360439, 42.45204917696383, 44.247010823546056, 45.96671691230397, 48.05491055502414, 50.14229286164541, 52.34026682960074, 54.35131448245696, 56.65810164943346, 59.33420868117409, 63.30477952981197, 65.9779105156523, 67.5126992984674, 68.8642530009826, 68.09050978821138, 68.04809583622122, 68.12102076328704, 66.13256924107944, 65.50801146097206, 67.52384081592413, 69.208309412895, 72.14993391151688, 72.40906169431895, 72.6653550917999, 72.88665041718045, 74.02533889434102, 75.82479322235575, 78.10240007906125, 79.8995591815051, 78.90256401682848, 79.96029544212969, 81.27399300238211, 84.06338781958013, 85.60023100901812, 86.68893384322307, 87.78004525527848, 88.86770805782278, 91.51166493220074, 96.58033630307044, 99.44268812544325, 104.30042055794954, 113.35719352387046, 128.86342236954496, 146.56405922690112, 161.40392384298096, 179.45447488425378, 203.6139564065132, 220.26569688881827, 229.25049380402353, 238.11940096531566, 246.17958004229294, 256.0091847713359, 265.0988408844332, 266.792095366725, 265.57266462033846, 262.13068482641194, 255.59685031043023, 252.8374876224222, 251.59970762002348, 251.85217434377435, NaN, NaN, 51.1317734690778, 35.18541565029005, 33.55568156807962, 33.84247547409337, 34.129276130928474, 35.15514818354177, 36.327709894272594, 37.49968337327512, 38.967744380796056, 39.98993210309952, 41.012837341209874, 42.183941478488855, 43.35353844244724, 44.966637715870085, 46.72599413566199, 48.33710907851832, 50.390939774571706, 52.59245877893337, 55.236444525534175, 57.58296987536917, 59.85701805803429, 61.76692489418739, 64.1612167679973, 66.73135781034082, 68.11988214067023, 69.18010794545731, 67.96608043870734, 66.0957618428516, 64.25203351298113, 64.44154227942073, 65.28420983075813, 66.59542958980929, 69.93517385429583, 72.94717834468014, 73.8592478092067, 73.04931248921379, 72.97312461129154, 74.66044670742902, 76.19502752343347, 77.58433347287874, 79.23271505808647, 81.43227286984636, 82.08579588967633, 83.83878393198502, 86.0345168913596, 86.90691987883751, 87.7720017536275, 89.5243265075933, 93.04528688528714, 94.79736032216337, 97.44741165377378, 102.7479710546618, 110.91870590457589, 121.52433980236779, 133.24665836757336, 150.76090816118753, 169.86137399279963, 193.31984318918705, 212.32832127159506, 222.9025578498131, 234.1681757983189, 244.8843161025506, 250.25082539185522, 256.72889732700895, 260.8674731944062, 264.84356468880134, 264.49444821915654, 256.8311509379599, 254.0435440703565, 252.0588437017123, 251.9915140436925, NaN, NaN, 34.262879074662706, 32.634840261705335, 32.99873413082677, 33.58152876554952, 34.0889171552317, 34.966026195543975, 36.28552680598321, 37.19781105228635, 38.18371496213357, 39.17033086902794, 40.52584366461859, 41.917966597706325, 43.9376031945736, 45.3640982003088, 47.12281237451112, 49.21401726615635, 51.413391201133976, 53.46605283867503, 55.22179343712757, 56.50193840938636, 56.49664742648443, 58.994225884809445, 58.62325988176222, 57.44468277398659, 59.72076670920724, 61.26629318224823, 62.58013724075413, 63.90752660543854, 64.1995393432148, 63.98007736353169, 65.66727976730911, 72.50411728460527, 75.22509731715753, 76.3347719291531, 75.22394807091786, 74.04248187676001, 76.0319000399295, 78.45567109430415, 79.84187177895353, 80.57012927256052, 80.78020867483043, 82.79503677098674, 84.06661966168299, 83.13785390871318, 85.14723791905192, 87.70447595799264, 90.26888084876519, 92.83272990898523, 94.47319159297162, 96.30702754480168, 100.16992227525475, 108.07475204072003, 119.13400007750474, 128.53154455213084, 145.72041548435033, 168.68605877896505, 190.0265902494059, 207.19671568300652, 219.5719738598131, 228.81614162940375, 239.20566281022124, 247.7521440634587, 253.73582960664862, 256.3872976917702, 259.8825285240161, 267.5555817359507, 268.4117130288364, 267.6813282519468, 267.0502406982261, 262.8818442091029, 252.41071017337492, 247.60378085678587, 247.77432352765913, 247.96890946569792, NaN, NaN, 34.33852377103652, 32.52595127501537, 32.77759717283, 33.98756866543055, 35.23217142497529, 35.77563145494105, 35.438327452757996, 36.02031863030415, 37.66941526169175, 39.54080144844602, 42.36842660265105, 43.356731543840226, 45.815646075966995, 48.20291313355413, 51.3693065459967, 53.34854572109285, 55.07535676734086, 56.79932296082183, 57.85328822551961, 58.91330949540136, 60.31622295714637, 61.707836523889775, 63.69137585857366, 64.63985820195988, 64.56143059208539, 65.8128972307363, 71.5469558838277, 73.59519983513275, 74.47188281362942, 75.71798528832359, 76.67709595476249, 75.78918527010337, 76.08351639334938, 78.3605779614949, 79.16604086818779, 80.18056251843268, 81.49481847464101, 82.06945316010267, 83.01407260439399, 86.38436207467096, 88.3527557466077, 90.5535369976915, 91.6437831270014, 93.64818097326888, 95.47809742595119, 101.17697718151335, 111.86532482888475, 127.17763364057251, 143.24344956778583, 159.13139660351658, 178.39297209458078, 197.9623654267403, 215.56536602544654, 227.387203688999, 233.79544470470145, 242.23330869889654, 246.40115473565092, 251.93204083691734, 260.94095283507534, 266.36108606180215, 267.4791169606709, 267.1619808264426, 265.27304300938545, 259.6228829714854, 252.33705688826925, 248.3926185703824, 248.3425618151838, 248.53574318892444, NaN, NaN, 36.739289887330884, 32.9711643945451, 33.40985692486786, 34.434979734917746, 35.68193903245394, 36.99995873515272, 38.058284333936854, 39.11841394599556, 40.32610313059294, 41.64688288898765, 42.78112569791842, 43.54492617942311, 44.752822202111616, 45.84871937705973, 47.28206652475435, 48.822590285754934, 51.06482465938983, 53.2641937036108, 55.539300426903786, 59.36152219202791, 61.34633298135983, 61.34039327130184, 63.027913017582215, 64.41138466844868, 66.0243686894151, 66.17020537424322, 68.01072312184597, 71.9157863829423, 75.5876302811044, 78.60382656041139, 78.82458241362912, 78.34028439173507, 76.5601151924476, 76.11492845466809, 76.8418336983604, 77.74542148123845, 79.31953961087825, 81.10896222342669, 83.37119994224072, 84.79560458761023, 86.87683368772846, 88.18833066868253, 91.04770579025211, 94.79228761157789, 96.32353811322079, 98.52013130841497, 106.47062711072624, 119.73475982367884, 133.9057856706273, 151.8599695235672, 169.3865365633006, 188.80254713959175, 214.43770015752406, 230.00382945233198, 240.88394144471803, 247.90819544071087, 254.8058696355194, 264.98866890360114, 266.87685425064564, 267.5025427066237, 267.57043272981224, 266.63910179730203, 262.2227376989662, 252.25050907538468, 248.36370026964892, 248.41612200464135, 248.71760783912006, NaN, NaN, 36.67058592712896, 30.169717571149484, 29.648865142845803, 30.968878781863776, 32.069258354898146, 33.53629625952673, 34.92713055006752, 36.612211610242106, 38.59326325136166, 39.46818147135966, 39.89979391309554, 41.586040677404, 43.64010358761106, 45.693374039067905, 46.933898593169204, 47.81330192641036, 48.689032329992564, 50.741438789378606, 53.16348735319967, 55.8812145808991, 58.11840436109902, 60.319303500879975, 61.93006220532172, 63.20916386464081, 66.13980308270045, 67.27892014038937, 68.27122224203072, 69.99175532015909, 70.83557188251947, 74.1063725665554, 73.62898242733154, 74.94982977517107, 77.59625729546241, 80.02538409431556, 80.68207157849739, 81.6651572301745, 80.96907317829319, 78.64863605267008, 80.1146509728737, 81.10416867826795, 82.82058338929883, 86.1947927512526, 86.92650116142387, 89.70856358031999, 92.93433392731914, 95.58451646517922, 98.08646237106278, 102.93629024067404, 111.63075908914209, 124.30662084862372, 138.03279991959855, 153.97909584353914, 168.76160065093396, 185.83046619985052, 201.2135228879662, 217.5728527448446, 232.84951242396914, 246.35897163420643, 252.8439966358014, 261.4231965811717, 265.8974765050644, 268.3772724173144, 267.4707964970133, 267.0891619457841, 264.91776450215946, 252.68187442565204, 247.94969671057711, 247.8031019406022, 248.20577718613006, NaN, NaN, 30.348742405552713, 28.16867061047757, 28.49511376358156, 29.41180575780752, 30.365681443946716, 31.31952728958485, 32.86063206668966, 33.85178414247405, 34.875734304257044, 36.74749241580549, 37.36529393585783, 37.945985217791545, 38.67624262879984, 40.14238102959593, 43.29825312723023, 46.162162930233876, 47.739649169555406, 48.87123320221508, 50.96229831297883, 52.320435267014176, 52.610056033324284, 53.379333952724394, 56.31073855882548, 59.61357967347791, 62.805329021021905, 66.47959358720176, 69.63147530002296, 72.82867848491034, 75.64417934323407, 76.44422108022933, 77.43102132790602, 80.1101297921342, 80.31833943876487, 80.83297141553861, 79.62737863621015, 80.91274652094741, 81.93478996634131, 80.76044940362307, 81.04675628358235, 80.276844354499, 79.61818567460695, 80.64291413112882, 82.6910756512115, 83.41864862290159, 83.7048732097865, 86.33720247964978, 88.97666491753913, 90.29499935803376, 93.23136715783842, 93.81272199088745, 97.33093924396762, 107.33120827089164, 115.86714316525664, 127.37882272954785, 144.50320929381996, 158.54080249311207, 176.01869989668086, 191.48337576353893, 204.11240197729623, 215.0879752390339, 225.8624805217543, 237.95987954675405, 247.80597139334282, 256.41148197158606, 261.8248168315665, 266.09435142799236, 266.9101197663576, 266.4441134221939, 261.75057584741637, 254.06707062847192, 249.89647052752372, 247.95026927207988, NaN, NaN, 29.950680886926456, 28.656483008397075, 29.316028281744465, 31.117844054769694, 32.25499349223071, 33.611713890642065, 34.450182464281056, 35.144497934129305, 35.72870855795814, 36.313307617928245, 36.491474972578956, 37.84533757902916, 39.68107531279759, 41.585750678828575, 44.48779623491082, 47.27813938644725, 48.85165916019006, 49.68845587101894, 49.86696112633735, 52.58361219501801, 58.05942311839072, 64.44839132735899, 65.17974331943888, 66.05227755306977, 68.7660772080461, 71.92845427020177, 73.98861639879776, 78.61924720596129, 81.2593018273514, 83.16985232115803, 85.43675611537032, 85.36394286766183, 83.30166737749391, 81.97284863869706, 81.67525314283674, 82.7796482954842, 83.65542801118195, 85.11504690311594, 89.37655027122246, 89.8087222893382, 90.82842224934012, 92.43413387311165, 93.45482967417193, 100.65240706030663, 107.58442006677815, 116.13961707088313, 133.87812337851727, 147.0114019696071, 160.16607400386235, 174.38183016003666, 190.72418902875572, 204.11762794484207, 215.82449389135562, 230.57534540432545, 236.76971604938484, 246.17108952343614, 253.74294064928796, 259.3507183593953, 262.9493737691629, 264.63184397158983, 265.33353884758566, 264.0817823979605, 259.13684589882183, 257.1473870935725, 253.17749489218863, 248.54533222348886, 248.13997785617204, NaN, NaN, 32.89493370169752, 30.567843587599715, 29.64292213467525, 30.338383412801637, 31.65893578892389, 32.870202289030885, 34.006941640233535, 35.03293423658797, 36.42574133354608, 37.194863647011566, 37.88613271921641, 38.98456837550121, 40.48536021235354, 42.872481146437664, 45.92235312775038, 47.64249282048605, 48.22100714391904, 49.42527285209523, 50.44689166694869, 52.0571591210003, 53.92649517340292, 56.20125776304252, 58.175439251383935, 61.18169709033727, 63.22707049134655, 65.57110670021642, 67.69598693628129, 68.79337550968995, 70.47580071653341, 72.75086586531654, 75.25152441745118, 80.4662190891116, 82.51556066999918, 85.45780441040893, 87.00054672212906, 86.41513418402488, 89.7164576265294, 92.42544853195982, 93.89107202659078, 93.23611803502268, 93.63828372760025, 96.3927655871533, 94.18685383099955, 100.2409304254491, 100.79991607822963, 105.57018674478344, 115.49873087616729, 123.97412887954133, 137.2856613050069, 159.49971862897212, 178.7731251364426, 198.16682811986087, 214.04837059219776, 224.8919945886474, 233.38139144348062, 243.64404597652688, 251.70981430774296, 256.6575639178689, 259.0495477615819, 260.0723247187183, 264.5428928118693, 266.5111122339867, 264.5443452737095, 259.12531423721254, 251.61564935286373, 250.33244513474955, 249.01783831480768, 248.845203055696, NaN, NaN, 34.77472301319023, 30.272019882596922, 29.901824250395574, 30.634915173086036, 32.547929593951174, 33.86597675229869, 34.8923072139076, 36.91553137378167, 37.71733126413065, 38.41086428040415, 39.58515131020383, 40.6853562989706, 43.365391022895984, 46.07998506055057, 48.684643692528944, 51.66189543078722, 55.18770416394941, 56.17232075180884, 57.05156122687263, 59.98836662819903, 63.44491136165922, 65.42012562513716, 66.8880372031426, 69.97132553302069, 71.2838707649608, 72.16499845108068, 73.99744854177084, 76.27092441411234, 77.58919034412857, 82.06252673043807, 84.3465019557922, 91.41116642133166, 94.49645248159601, 93.75881811213745, 95.81236149492942, 99.47393368311516, 102.55439863830814, 102.62387699756373, 102.47727365186824, 104.02325442469089, 104.12986926383657, 105.04883199491877, 106.69672596256804, 109.45727945772269, 114.41918907426218, 121.4063396492537, 128.77986792187352, 138.36520243758994, 155.04704806639106, 173.94265212054557, 189.33021208583747, 201.80069923827807, 210.56454824388436, 225.0682733461202, 240.5928914916674, 248.2921450922541, 251.95613069968184, 256.8081452145644, 260.69043489675664, 265.2796866647047, 267.3972280906039, 264.76071261044336, 256.30089739432566, 252.2280645121218, 250.84638847943867, 250.30760935010892, 249.82260472708722, NaN, NaN, 28.204419183048643, 28.27598739182182, 29.452734777326796, 31.291426420886726, 33.42515454582815, 35.48244526873472, 36.359024527925655, 37.08803354497802, 37.078110450568225, 36.85392430739635, 37.06920768686347, 38.39004195597616, 39.70981578998093, 40.733208462944056, 42.71373992186032, 44.32734082655062, 46.89720010211287, 52.484954512403235, 54.984572227614855, 59.4632407734596, 62.62376837866473, 66.15502321405455, 69.01499642061654, 70.99879867067135, 73.63408255457765, 73.25962530330015, 73.09803885884035, 73.82877599227184, 76.31361336965891, 77.70743625595838, 80.64146613308428, 82.76130254302167, 82.90185733777048, 89.14319100031024, 92.90198517696105, 90.10195247116279, 94.65985607879992, 98.99868680062077, 98.20063330769773, 100.02627155910547, 101.63864156059194, 102.18872341276479, 103.0919266723618, 106.21635952008303, 108.80314595124834, 113.22273997018715, 126.09235067820593, 134.9549844685848, 141.789497290711, 151.9598095025097, 167.909452306315, 187.79870428611068, 203.26988173232942, 220.0754496495025, 229.21434970538294, 233.6666020586287, 239.4066085320926, 247.7496023793832, 251.9482659720034, 256.6146826836982, 261.6285182787181, 268.76622665442704, 266.4260954562535, 261.7767198014735, 256.68376944581814, 251.31702547929697, 250.342126741569, 250.45093546750147, 250.78110053297607, 250.67505793013902, NaN, NaN, 29.344310585554112, 27.348923916121375, 28.156192673462638, 29.47629482568458, 31.09293306755753, 33.37128490211201, 35.72087741673162, 38.00108530998992, 38.58632894686018, 38.063639426457314, 37.687158889042124, 38.49131312791784, 39.21784898438918, 40.23822156619713, 41.40799515940624, 43.093847192056764, 43.97303060987014, 45.51126359277563, 48.665532206582455, 54.175412759485056, 53.54396997870787, 55.223466258433376, 56.98174541030652, 59.54943015962707, 63.94973825594138, 70.71012205985727, 74.37927338970194, 77.59745603342387, 80.75369584686615, 84.13470870027963, 87.51384431081064, 88.24129784322727, 90.36710238484243, 91.60834526587651, 89.90893736186443, 92.40121924915897, 100.11251862270458, 105.91516879621304, 106.21619206199863, 105.61653497213864, 101.82067779744422, 101.45855737620266, 106.42641902535215, 109.56670116599436, 111.2337370242519, 116.02179478675966, 125.06574387263079, 131.87856913959092, 140.58322008824965, 160.03383034683026, 177.58868438272032, 192.68294151308825, 208.32151893018505, 218.05207680641118, 229.71284929633458, 240.2141762784856, 244.83598963906215, 248.11122686456437, 254.13341249246167, 261.32799961214636, 257.77157181103297, 260.88250375093304, 262.0197502930601, 260.8803904524508, 254.71780255927516, 250.70726448798084, 250.08647422396388, 250.4087831205672, NaN, NaN, 30.91089524319357, 29.39467423582652, 30.829210910548763, 32.22554592400043, 33.4022059748084, 35.38663550722963, 36.930597166194126, 38.39731446553491, 39.12730603507649, 39.967050087414975, 40.80644483992301, 42.12532723688825, 44.14030675058558, 46.34243818215392, 49.424333648155084, 50.33705640216491, 52.5756555244249, 53.41630390527763, 54.14861638051368, 55.20760509154346, 57.11570912096584, 57.842750198341776, 62.321588203517884, 68.55601090018031, 67.95690467574033, 70.88901894096533, 75.80862391362787, 80.58149609300023, 83.88552270753833, 86.89276154316897, 87.70435313276342, 90.19582271418588, 90.41801536836293, 90.05020854509316, 93.1315526575578, 97.23090710114406, 101.34283707570648, 104.94434697015551, 109.42549360941622, 112.50262146393328, 111.37529739266108, 115.79530164611721, 112.14627366351212, 119.15077774809066, 127.64478544851961, 136.32416793021227, 144.6212020810981, 165.7283989422765, 180.7315112245882, 191.85685382354933, 201.62585088984827, 221.41623861003336, 233.09322834513597, 239.58284814622476, 246.18312867700652, 253.38916397011442, 258.6589197371901, 261.45806823653237, 261.9314283919187, 264.62431481495884, 266.2599919530258, 267.2490140753673, 258.3041926817653, 251.26626387476253, 250.58946243806267, 251.10078631093364, 251.39407686286853, NaN, NaN, 29.3906830017219, 28.280025765599678, 28.49729242458693, 28.714217343946363, 30.1105920949601, 31.615961831044498, 33.04846552738428, 33.89249483890869, 34.847237832026615, 36.94472149860481, 38.77943267006252, 40.39168548557354, 41.01097266915071, 41.924040855272075, 42.79863609496476, 44.89231124853754, 45.94646257785686, 47.85409241641305, 48.58080229282667, 48.099473863307345, 52.688479142949156, 59.23199426555484, 59.88647341429239, 59.14360786496564, 58.767387390995616, 59.78848276187809, 59.710534736519755, 64.9227723137807, 67.3467604404159, 70.5740254934724, 76.88578783318684, 81.51063293951152, 84.79973904929712, 85.73663916969367, 89.99338744653966, 90.50810557172152, 90.72745325962966, 90.21327127273852, 93.52253274595404, 94.39421230401078, 98.11066324532074, 104.37583339288153, 110.0695994103557, 112.99788239808407, 111.35972247414584, 109.71802204807186, 116.18161653494305, 124.13582721187028, 135.95573953308718, 142.21428092988157, 153.70808809547157, 173.65641403056708, 180.9146016542522, 193.33129160201526, 214.42266319948504, 229.7381563564433, 234.654874126723, 236.75755905625957, 243.67926407754194, 254.97375937300134, 255.8098796542776, 259.67219942647233, 261.8867351499456, 263.1155846831427, 264.81379423731215, 266.2598617862924, 267.67596786368244, 262.50289995939346, 254.21874940899406, 252.16407318639202, 252.0682268892406, 252.39565580978652, NaN, NaN, 27.065057154124446, 26.764161716415213, 27.53481026537697, 27.603354024626167, 28.186082188886616, 29.69376534786583, 31.456169413742497, 33.182279157244835, 34.94562851171694, 36.488794800676594, 38.14329686985148, 40.421461287234926, 41.48260204881406, 41.880820321116644, 42.72006006738944, 43.85404977921425, 45.249617674872844, 48.517992668665435, 51.967705724700004, 54.4992756789453, 55.85122061427953, 57.535328912538574, 58.93155210616161, 61.20858931044499, 66.93933170755841, 73.63180105893746, 78.76584797262876, 80.95996172535332, 82.79189968305184, 85.27613877185833, 90.33367766361295, 94.80245240693039, 93.4117062233599, 92.02269916365785, 90.98400954163878, 92.29703931631684, 95.68428224207055, 102.30677100938308, 105.08167265397293, 104.34020350033039, 108.91526303432745, 111.56580067687672, 111.80904192540898, 121.13290675423495, 131.77239578506888, 141.0903488595326, 149.7001980579794, 168.7773963412649, 182.60356472830745, 195.5148099059472, 219.67671722138306, 229.54342373106448, 235.8968110019359, 249.7491088981033, 256.65678829121947, 259.78642447876166, 260.77335521300233, 260.8119620812434, 261.594666040069, 264.37179382163794, 266.3952337993557, 268.40573285411796, 267.0226877180711, 257.96759876814787, 254.9543642869718, 254.92369969984446, 254.99616382555627, 255.1723251547375, 255.37685082345575, NaN, NaN, 25.3746197408656, 24.337985360511706, 24.88613171592938, 26.0234369248167, 27.602985722048494, 28.44393634046211, 30.613471202091265, 33.00411097742049, 35.69055795100971, 37.56324827780582, 38.6990719509699, 40.05685656418298, 40.74982011318011, 41.66274354805312, 42.168270262087404, 43.00567191263895, 44.32367573776685, 45.34920072204572, 46.260518339014205, 47.87006531216568, 51.46876816375695, 53.89188109124194, 55.209255219537184, 57.51637230675087, 61.373351474109036, 62.68440576245977, 64.32656637260457, 67.18427322241173, 71.03497468876881, 75.9998160599481, 80.40474856817941, 82.3805544624006, 85.13566299924584, 88.55703422561756, 98.58472888931105, 99.46681508652003, 96.26557865894937, 107.83991640789716, 112.92827642152552, 113.3821697826291, 111.9281824658814, 111.95041548865085, 120.39433004851124, 137.5350095641768, 148.47004473515938, 156.46169729929483, 166.45793158076546, 172.39471056572995, 178.28410854259675, 197.5029919195193, 220.14843416811877, 231.05747817297376, 244.59000787112905, 256.67914451718536, 259.07645505372443, 260.0551232097085, 260.69406010685765, 261.7434305625877, 264.1195236081656, 264.14709042244874, 260.4163140595703, 255.97299690192594, 252.4582354809795, 252.40712552575002, 252.72833831894914, 252.97818727770326, 253.0756772961405, 252.97192652561867, NaN, NaN, 28.02142162214453, 25.991229061872893, 27.60648273812048, 27.89546536687357, 27.484290479867813, 28.61835739777716, 30.306608237205044, 34.05885035173562, 37.95603912878472, 40.4520605725567, 40.9598985309769, 42.13306981962367, 45.43704370846285, 47.82406628495125, 45.46581057664579, 44.941387916401794, 46.40593585159415, 47.97876282053871, 48.815968739556205, 48.953695498363885, 50.932457485813885, 54.35278744752852, 56.56143061717877, 59.749951787009, 62.82712257244782, 64.46804950532055, 66.55131200142834, 69.85173504547573, 73.48260740259953, 79.75944978606914, 81.51907960838646, 83.940532659968, 87.24774458612369, 89.78231179850103, 97.59356701193651, 104.65373386244303, 117.10408470263928, 117.77936525480021, 113.92026321926046, 112.60915531326758, 110.58435796726967, 110.61557396432214, 116.81771954858566, 131.8394529907877, 143.17358273230022, 150.3566897654903, 162.2067962663, 175.80293540681532, 201.5187614902775, 213.40131337852347, 224.60617411555526, 231.74793477415872, 241.2675121301503, 245.14421214685657, 250.22463892675506, 257.9349207674198, 260.7384242465362, 263.3976798262921, 262.2876066410975, 262.18798465330224, 264.0262897780342, 264.5140541788742, 264.9556291948502, 260.5636027753833, 255.98286299461506, 251.19611675481218, 250.28068770645075, 250.6059703313501, 250.71804975182255, 250.9746080078453, 251.08881536934578, NaN, NaN, 26.76856750016089, 25.32877648974365, 25.80309366553421, 26.90357863395794, 29.955673304339175, 32.60614515004919, 33.70591759472315, 35.06421896555176, 36.273204673489225, 37.48367025040769, 39.765009020890304, 42.07794761153275, 44.94014680337327, 47.843322590721066, 51.480115348012006, 52.90732072198371, 54.29195921243125, 54.50302963106752, 54.720088671912265, 53.72377946646015, 55.59283255251073, 56.134239119671186, 59.21035051682415, 59.75475684278233, 59.302735414161056, 63.925713570626336, 68.98811504352943, 70.4132547665286, 71.94676223977565, 80.86127902539634, 85.92368543586042, 87.0381766295346, 93.54463243552011, 103.12053483781668, 103.45526094726924, 101.90548165514365, 102.90375763604625, 103.69537911732408, 105.13775476409144, 111.19772451872194, 116.69832198670993, 122.4558401811945, 130.8477796499813, 138.60906700523208, 141.06887235280945, 139.30602342447065, 152.91177509020892, 177.88224201762176, 206.06277286846756, 220.3386216263845, 226.86255170427182, 231.51726522146484, 238.74137101036985, 245.1702987267106, 251.59923085717526, 260.5906692459555, 262.8232644911844, 263.99487283218326, 264.7135661460247, 264.1145198261076, 263.3405739567716, 259.91054490280555, 257.29026308107194, 251.6050525532619, 248.23752266021106, 248.26364541432352, 248.5177914604486, 248.76702837247973, NaN, NaN, 25.775838582447797, 25.73558943323872, 26.544582152314067, 27.867550257837856, 28.821212286585563, 30.141300487549717, 31.277027296368615, 32.37657618264209, 34.13881202165719, 36.6015378527773, 38.582402321290765, 40.48675157979866, 43.166841029201116, 46.07136965091851, 48.42033290579584, 49.809693739971735, 51.78618388399232, 54.46668153867915, 56.33843046616094, 58.28454198551016, 63.788949522649546, 64.22344054790823, 65.65164805604516, 67.95552289366488, 69.59622543316587, 71.4569380735104, 75.42576228733073, 79.06025436385809, 82.46674737681798, 87.08991377481284, 88.2949907144124, 89.17092138171547, 88.50498535127096, 89.71039492194663, 93.78892417539534, 96.44032455070942, 96.90233056724603, 101.77420808370559, 111.91150569022629, 115.01434055834652, 123.77464342959125, 131.52156460144028, 138.24538279979348, 143.93953277711233, 141.35148993152384, 149.69906015059135, 167.68962637548705, 195.7720918208695, 213.52619151059122, 225.9049738467965, 234.97905331167965, 239.0085740329833, 244.77832576454898, 251.48964225500842, 260.6855886772097, 261.48686563619316, 263.1385954142184, 263.11062110534664, 263.9749828599073, 258.28105917842475, 256.5890045224235, 255.94585518040765, 249.5097169180364, 247.98752533673365, 248.24322659502317, 248.2741685910718, 248.51761556154761, 248.53405637128583, NaN, NaN, 27.475356939913123, 26.843791135871673, 27.61304060131686, 28.381638448972293, 29.36994348792098, 31.13404794597969, 31.829234631244773, 33.554080741630344, 34.50892167123228, 36.6727489061427, 38.32374340121133, 40.451323082479725, 43.35037867934392, 44.268895598124786, 45.69461463755858, 45.86937178586535, 48.77210403803316, 53.075300336481504, 56.67501732398095, 59.46147913740105, 62.32212317286818, 65.1831134769405, 69.14657940417999, 71.89604858876686, 76.18678890063346, 79.1582766124879, 83.0105487464516, 85.20838714403187, 87.51616083018342, 88.05103465756704, 86.07341391986547, 88.49658343206346, 93.54793611227068, 91.44243804204599, 91.54743838385974, 93.41580515363205, 93.6335144978924, 92.19590069214057, 90.76959668674132, 102.23133799140284, 115.12312270970473, 122.8614273098745, 121.56268407778904, 126.89551041433704, 132.88064643811603, 137.76947185323127, 150.4105110443259, 161.07932032463037, 166.39112018647234, 169.55637112695095, 183.24143473334036, 209.4602151059541, 227.22909179557803, 235.4994249412514, 242.17860529362778, 252.4151515536774, 260.0275060830699, 262.002822840847, 261.9801843753621, 262.984762376922, 264.51763556077793, 265.79667235561345, 265.6353503783549, 262.5867971650239, 256.8529704491016, 254.93551060751534, 251.57033953195304, 248.11167287404527, 247.9991656515376, 248.17705815648546, 248.34892685984227, 248.43835960514843, 248.62468367976257, NaN, NaN, 25.47713216015721, 25.068868023933923, 25.72853848101566, 27.972932316784966, 29.738564604229186, 30.579119559636954, 31.60483925375729, 33.88429794797032, 35.090764636047744, 36.22764694108948, 37.83944540049761, 39.59827045498865, 41.57405176893084, 43.00257955046995, 45.279839384408646, 47.95840046221004, 50.30767036050717, 53.35632869407, 57.02882626835944, 59.601300222274354, 61.24662171854408, 63.14387861285935, 66.66400788987737, 68.11755825625013, 70.6085344580198, 74.42549694140696, 79.25918625288399, 79.54142613607077, 80.55720437002371, 86.57517661279088, 91.56738545428618, 92.15063633110316, 94.04850582787941, 91.26655729537323, 95.37342952131306, 109.31953309867498, 115.34033238798563, 120.9467100305031, 127.42423550291015, 137.06356736273298, 146.3081366637691, 155.34280683736532, 159.51303303223094, 157.83527229091618, 162.77834847070656, 177.6529038468996, 192.55300334217785, 201.70520996702996, 218.07029875112303, 235.04747732101407, 244.563205529786, 252.28490969191733, 261.25526188125093, 263.8416014151932, 264.25507055440477, 263.6459344875968, 265.7914295153785, 263.8762267436324, 256.4247499380388, 250.62732217189648, 248.0806772477884, 248.06803981279342, 248.28633962219186, 248.3889293689058, 248.52382083343971, 248.5815921911626, NaN, NaN, 27.4413371438828, 27.29085241702471, 27.508278002490496, 28.314516827106278, 29.96833618381884, 31.364974176463704, 33.35103469084179, 35.039621823508995, 37.869442464798816, 39.59230695837892, 41.16962664216967, 43.044560294895824, 44.88693069506303, 47.382443069412446, 51.90532214204061, 53.73828067290166, 56.011395717315416, 56.14995903148249, 56.65952359973792, 58.7874823047104, 62.71071648698952, 65.78783052834646, 68.53549114330218, 72.83145328054114, 75.0252363483373, 71.70635131264532, 68.17283623618872, 76.09621215031784, 81.49121545794027, 75.54630545673328, 76.97059366964, 81.03230587465927, 93.68684542412106, 102.71322501637309, 106.5735471267478, 110.32434940932197, 112.95832941449798, 114.93544973247604, 117.23678060001568, 121.98309221618445, 127.4179711339016, 135.98617692606166, 145.63209815463165, 153.78546375743292, 157.7802931297863, 168.16531366519462, 171.2561591815013, 173.64852086934056, 183.321984987941, 197.47015308582246, 211.6091200962555, 225.94200419111763, 239.3644792910658, 249.17334856554402, 254.47339070393787, 258.600071920737, 262.27110995300313, 264.4189542781736, 260.5566983655248, 256.573073824126, 250.17900237443516, 248.1571640118478, 248.36654689095533, 248.6570969983526, 248.82930075482616, 248.93143126800803, 248.9957861110171, 249.14832676081443, 249.26554137447485, NaN, NaN, 25.29193043587565, 25.436276566570783, 25.839207969638764, 26.387500457127636, 27.414203509934488, 28.369615375381372, 28.91633965644689, 29.8303301887229, 30.7096251626227, 32.288517519926096, 34.38442784078538, 37.43721831908197, 40.11727910404117, 44.161747443311114, 45.07614749710063, 45.552837524193734, 48.19494093419436, 51.76229767026951, 54.07832059504658, 55.43744857313853, 56.7968500247552, 58.921379345384324, 67.22293745821005, 71.33844890500477, 71.33337911063202, 64.93703592253078, 65.51576360598906, 67.7130615779665, 73.43652099217144, 77.62388020258528, 78.12574210794811, 80.53932701550595, 88.30418745997734, 96.3854814167237, 98.72294164438246, 101.79429581008877, 105.3230218090069, 108.62408480791376, 112.08587903878866, 115.91280188599981, 119.80064710870562, 126.7197315406321, 132.75741026037656, 140.7432801431691, 149.64026187892264, 159.4049913219207, 165.79410954296776, 170.54424024340946, 177.24163859412366, 179.75105755810011, 189.36117378502107, 196.9602034532241, 209.38557671128208, 226.378126647599, 240.59925093082458, 247.04416365448316, 252.75732487317785, 256.7673224769038, 261.40842765813534, 263.07668813668374, 261.0630511462874, 257.33970975859097, 252.5604880367636, 248.9595647417571, 248.56989340229984, 248.81617224645868, 249.00033685422287, 249.32748157572175, 249.35225485503491, 249.44397426660242, 249.61957761227308, 249.43861886136702, NaN, NaN, 26.54787631132624, 26.10201733820591, 26.61363860360701, 27.050433351026058, 26.973010505325515, 27.04203207659611, 28.58407439482271, 30.794764965581344, 32.92687010283123, 34.76216932681901, 36.964702470692615, 38.42828168121387, 40.85004810721311, 43.644565045073186, 44.234437836639025, 41.43305426641074, 43.26805931743352, 51.651107327222, 58.417065401953586, 59.739815726365975, 51.01643704743383, 46.665631922055624, 51.07120227974211, 56.87593932910791, 57.23830290096253, 61.13088176461704, 64.13360116399153, 68.89681390085107, 72.04618372304498, 72.11458735517166, 73.13000737666007, 75.39375875767051, 83.62220941774837, 91.03368527946618, 99.40085690791268, 105.35502859237249, 109.92557354918942, 115.37411724351887, 118.66869144158265, 121.46994935433206, 121.56075462659702, 125.98260596349165, 133.2639855929301, 144.73804492443463, 150.30355517763692, 158.0783346880274, 163.3737869349048, 173.9462911537061, 176.08164834819132, 186.81504982112992, 210.5854300754249, 215.97053631723446, 226.1780202753915, 233.21812451888755, 241.7979605565123, 250.24086008654328, 254.63762627147202, 260.13287932555625, 264.98273901647553, 265.9690585808068, 261.72414744018084, 257.5193584541691, 254.391028939696, 249.9061665589988, 249.2818561431462, 249.52185288097678, 249.8447385031828, 250.01469689375577, 250.10550668092816, 250.2130420384264, 250.33311938357713, NaN, NaN, 25.260580930295674, 24.81535723107449, 25.179344431967653, 26.2807043335477, 27.529522801910467, 29.809865672636352, 31.94122535328289, 33.62893003189261, 35.09836846113353, 35.97654069929478, 37.29934794425723, 36.41281568081115, 35.2290785776778, 37.8728863805472, 39.337559035856614, 39.99527774552196, 46.536840488856384, 55.139040533589366, 59.035826088668834, 51.83334402566457, 47.30185712595777, 45.38199762997657, 46.55068882998571, 48.45269929583195, 51.6763112061412, 56.078919165596254, 60.7868628542336, 62.69306613176841, 63.129205813425365, 63.71415446244231, 64.43645219204265, 64.4363013793461, 64.71736785385244, 70.8863558394049, 81.7649872892941, 97.48369653201986, 105.70759512705293, 108.3705189318722, 112.1981376374239, 120.12048687378616, 124.55619013653103, 128.76831044854438, 131.89812557889408, 140.0047434335552, 145.0018262639107, 145.8122464660295, 146.7631138725584, 154.30446684100562, 158.3853483806716, 166.37878376025753, 182.5128155206755, 203.12773442513102, 216.83198439199907, 225.76596908576826, 233.50446293558358, 240.599512966501, 246.660337059228, 254.2161160141926, 258.2984133326898, 262.1255068081129, 263.6283293988534, 265.77531654948103, 264.72558349906495, 258.28280926764387, 253.6826698611638, 249.2135900050899, 249.09287607674116, 249.34089265939082, 249.520273650807, 249.68927285610886, 249.86568516155276, 249.88443455189753, 249.92770902683836, NaN, NaN, 26.184071781814016, 25.810961311904787, 26.763665787521436, 28.45441536012877, 31.472335401932177, 32.12948481498033, 31.31557122741948, 31.458110710185554, 31.602387849563762, 32.04086772877239, 33.95245698942905, 37.77910944659805, 39.175708995173444, 43.36824214651903, 52.19620518380823, 56.24091636389677, 53.88783296645862, 48.58688464674295, 49.82860166696221, 55.192437221149724, 57.986880091646, 59.15468130358606, 59.00085597490061, 58.11945078968264, 60.17953290274318, 62.092785743613426, 61.79305542459421, 61.19635857926032, 62.069305711275256, 67.79834359132231, 69.99318519816931, 70.86696454175166, 81.7426018539226, 95.99753463636011, 98.33519059036395, 106.70853200540373, 108.03197621620306, 104.51020527642734, 100.09479472223677, 95.38932655041711, 93.436553307406, 93.21568378975992, 106.00866627727349, 121.89224670103843, 121.00153006498073, 121.21796095832795, 122.55635594334854, 123.67419285487017, 129.43130586456994, 138.5259418829157, 149.81842848362678, 167.16315230943601, 189.95265308158451, 216.06122852746282, 226.2725941656888, 233.34675839123992, 243.70789666166132, 250.06918074465457, 255.0192728662893, 260.1453931398989, 264.47865430045596, 266.39332709070743, 262.8722330362167, 254.5932315767152, 248.81158531251006, 248.348445407045, 248.67638044621484, 248.91995320178188, 249.09249936523136, 249.18796099383138, 249.28028662799835, 249.3748714717579, 249.42195402585298, NaN, NaN, 26.375201842524017, 26.963553715954408, 26.88669313965762, 28.430432640362977, 30.12243298330537, 30.707892639130584, 32.54668843894411, 36.37077557111482, 38.205020315283065, 41.29667959182936, 43.64937169797108, 47.03202036320535, 52.10265844522008, 55.55868240784596, 50.10949812472293, 48.03444922088364, 48.02367145770331, 49.044738658750425, 52.49934402383948, 56.471785700838225, 57.06197881500344, 58.382766326703404, 62.796321609909846, 70.18044103754343, 72.38372355688765, 65.2049157225826, 63.322445775538036, 65.74325857506305, 78.30611238966402, 91.09547835924171, 99.70188644697109, 95.86473269350714, 93.66631871231316, 90.78864556199558, 92.98471732989431, 98.60217813064777, 103.56729087754377, 105.88613128139389, 110.29357593656506, 112.7055767922831, 115.05672239877003, 117.39045415670054, 121.26881733568028, 124.87199825441367, 130.5675171137305, 141.94503566632665, 159.81769104848664, 179.8874327877044, 210.1058513081076, 223.67639017702683, 229.4930466480635, 232.90756545001702, 239.35913265755897, 245.45202391889492, 248.6568150105624, 254.91643880157824, 259.5314266056044, 264.5234397118514, 265.5758554268032, 259.10955615704484, 250.65616118179167, 248.26113138562155, 248.54331903981637, 248.78583125722295, 248.995431644047, 249.1379655294313, 249.2329787319012, 249.3010602209048, NaN, NaN, 28.524624760945606, 27.48660266823192, 27.702253080621276, 27.40175716386555, 28.871914136781605, 30.34003395138896, 32.76575449795707, 38.44065478363825, 42.045321773091814, 43.73255702081046, 46.080173970922985, 52.18738499325232, 54.16161583010626, 50.483428341476376, 47.82162576900876, 46.930093408636694, 47.28524363834449, 49.85336972537146, 53.969732645946884, 60.515631860199015, 60.77212543970899, 57.12196699641258, 66.60384060885269, 70.4694832336477, 64.9473074337667, 64.827706790094, 68.0140847182008, 72.41430374515141, 80.01826430865124, 89.3822451800162, 95.99269441571745, 96.99230947128926, 89.82359587256022, 89.71914208591919, 91.37580779244716, 89.92564784659959, 91.45339580479683, 100.05646686964103, 103.36503427176937, 106.11514447631004, 110.51439823233285, 112.93715013988793, 115.36741992759805, 119.36406828483975, 121.35847543974371, 129.35949295153534, 152.91247713864277, 170.2804004931087, 181.15802087820393, 194.06133331110146, 213.93572496365383, 225.9111767353512, 232.24559225156688, 239.27614354319613, 243.90720752900822, 251.2322750162173, 255.58490870225913, 259.0880441781199, 262.4028311656509, 264.77728029721624, 260.10604490679077, 250.31526602777848, 248.74121306429646, 248.90816900872565, 249.30235627939223, 249.36984127756907, 249.42874650863115, 249.49826889353932, NaN, NaN, 25.336733036364762, 26.88304468835589, 30.202427173981945, 27.917256211418334, 27.17239715180237, 27.45955114087259, 28.632590393657082, 32.31347604814368, 36.36082242925942, 40.18761279127388, 42.391070880237606, 45.84684493459398, 50.40040436835477, 55.83583052347555, 55.61206972656554, 48.40124988715214, 46.844759863161, 48.38040544366545, 50.50850253089235, 53.515249162792635, 55.16627642205707, 57.14644353299297, 57.2147713769451, 54.78287880004645, 59.77634957897204, 68.30395868726433, 66.53281367610255, 66.2273115881106, 71.43568302532744, 79.36780334015259, 87.81932267092077, 94.21608957951703, 93.4866863893261, 87.24027942758134, 87.02133291677465, 89.3734049893825, 90.39364987336643, 95.01517679273145, 102.50439983624412, 105.2336655313307, 109.32155793052799, 112.64192924163132, 116.17291627260033, 119.92233350580872, 120.35981978536094, 114.39720985850448, 125.25403316777482, 150.31984351777285, 172.36839551723867, 196.40529580709, 215.8113187841019, 227.17147424927686, 237.86004536841432, 242.50719180524396, 250.79356957297384, 256.9581740950406, 261.8373435727712, 264.50707949899373, 264.3173751165219, 263.6642380667257, 254.74471816243727, 250.0458915660735, 250.20686258724405, 250.52376584661528, 250.7612750612045, 250.8623558905093, 250.959230459194, 251.08014601835407, NaN, NaN, 26.14502415683362, 26.657711574765862, 29.752702302648885, 29.60548843910195, 27.390873628957607, 27.16245473505795, 27.893212693433753, 29.656244730509023, 32.81971393577872, 35.90781321230436, 39.66033240022343, 42.60253635060912, 47.67881466895665, 53.12111226420879, 52.3211233494489, 48.48408159741287, 47.51479188928648, 49.124867648823674, 50.587091898627605, 49.845865024289886, 49.32775553198909, 54.479188248721556, 57.0498268663009, 58.435820947835396, 66.73976993424256, 66.37357977997952, 67.16934090719279, 71.05922749924743, 73.2584856977764, 74.06032517419645, 79.93307543550104, 88.38844144369854, 86.552341587527, 80.15036456904924, 83.97883634694253, 87.94393680775791, 90.06087118947528, 93.07172545737284, 99.25272416076699, 101.82836158462896, 110.14040850313968, 111.02786115071471, 111.90037474630087, 115.85731352386847, 117.60408747820969, 118.47320907923566, 116.92810888818957, 111.64270002867462, 126.88011660087814, 151.30459835240592, 171.78881934859172, 198.52484004472768, 220.93948426161728, 234.80606526953878, 242.56837257125028, 248.5779982329011, 254.03742065371654, 258.461095594825, 262.70866453278404, 264.76280519270153, 265.17818750360607, 264.84278210750006, 260.81717471550775, 254.62160798932123, 250.12585944229247, 249.78485248481402, 249.81618818169298, 250.0535367588493, 250.16713020255213, NaN, NaN, 26.142538464020042, 25.62218999699626, 26.505915524501763, 29.597243164215673, 29.521501790607118, 27.454544929926367, 27.74382220757325, 29.581351314553633, 31.85773833586154, 36.27289502673607, 40.02472830449859, 42.375602391323945, 45.31647872976131, 53.41340699721835, 49.74111560160931, 47.67262393901346, 48.77077505230584, 49.871082316487914, 47.66378739470989, 49.134781033533365, 52.92409066661417, 56.818593501845875, 56.22297358642148, 63.28006885572088, 69.52374135242556, 69.7383597199135, 71.64219864705395, 71.27253695510376, 75.09253092448044, 76.20010031529974, 78.83616471988418, 79.57120516387481, 85.01528197435414, 87.43859442209276, 88.1517608772346, 89.09308081026293, 94.31197628572151, 99.7456014128999, 101.66319469555765, 106.95805673412802, 109.9008539873766, 110.12107491355503, 113.86275413830084, 116.93821434890349, 117.80550518272719, 114.49971237688641, 111.41791422137089, 130.44728936724155, 150.88891631309997, 168.25854773473503, 194.97189234544615, 214.79629314531965, 226.53983179988725, 230.52956258081926, 235.1408189915653, 244.4362810425255, 251.5138608000158, 254.68642655939357, 257.19554611494596, 260.99745546526395, 264.29371876754635, 264.50968006584816, 264.1224443073898, 263.7315433605716, 263.13715025826957, 258.771499391488, 252.5178949068316, 251.73956389881863, 251.56954251949125, 251.8893595395542, 251.93386672544023, NaN, NaN, 27.656462841558803, 28.31567584523367, 28.97477983089107, 29.707865840869864, 29.559160000574725, 31.471070471035286, 30.29001427813427, 30.062101695789405, 30.42093782404515, 32.69829732930233, 36.07857629919399, 38.13135708219461, 42.17981214374995, 44.7524966366233, 53.21278700931112, 52.85670018554499, 49.39082881064332, 50.341998820396235, 49.38256849208505, 48.11912600092063, 47.70485832980972, 51.523508771966156, 54.24244052871618, 57.69430404771514, 60.417044448510815, 66.14713308771444, 69.52346015296945, 71.35073978076942, 71.19249754653104, 70.08400847670427, 78.45479544102274, 82.78870305392627, 79.62665444633329, 83.3770161691193, 86.682064344557, 88.95273572835433, 92.47739801190887, 97.92314240621569, 105.78950752834632, 111.45414754459219, 112.71234829482303, 113.8083178645885, 115.34229147817709, 116.21425597953956, 113.3464697691129, 114.89494585388088, 124.61147774351998, 144.10267961779533, 158.8054812914272, 174.16243197007338, 201.04567975284263, 216.72384047283376, 219.62584315464477, 227.16893502817044, 242.908603214535, 249.97496002983095, 253.24124418696772, 257.5760981165106, 261.1978847645595, 263.2057363158796, 263.4658283107993, 263.3880770843726, 262.7969876396087, 257.91482918027145, 252.74494720514355, 251.82016236645126, 251.98231239636021, 252.32581890436117, NaN, NaN, 24.22607693110948, 25.18196075200939, 26.726476097875043, 26.35485306840534, 27.08922911644757, 28.929097575432255, 30.691727788409946, 30.026937582921477, 31.793006193928747, 34.8069366757992, 40.919484858039816, 43.34162969722423, 43.92038646323408, 45.16705899597697, 52.07981210558212, 59.28942491126813, 56.785871026120496, 51.40516140650765, 49.780977379893635, 49.47912726797981, 49.91428635872989, 52.33500470723772, 54.544000085634785, 56.85852888570666, 58.068383901067804, 59.612173852234285, 64.13275628781811, 70.7491361877595, 73.50364829790888, 71.72835867496876, 77.8925654645289, 89.12694670169252, 98.83563816556507, 87.48775641942566, 87.82229666299114, 88.13445402176636, 88.11715016979714, 89.6485078217044, 94.72771285855409, 102.68077953935374, 108.90382489935264, 113.66717545521065, 119.16634901765016, 118.9865982065788, 119.71666767587045, 120.63613141613402, 125.07108589431263, 134.1010467423847, 145.58093023378814, 161.53990560112973, 183.13687248940843, 205.41060571979003, 213.9735385072775, 215.4098669133659, 222.35102348732414, 235.40667067417624, 246.075623967136, 252.06452179151722, 257.6644030907056, 262.1460218544027, 263.99010509364643, 264.1682216738475, 264.0680863902612, 263.449823808586, 259.8717177565699, 253.3373643995916, 252.3460135905204, 252.66481733506677, 252.76528928056277, 253.18096355434417, NaN, NaN, 26.853028010899482, 27.291414603041368, 27.50978652321319, 29.71570440130117, 31.698235378127084, 32.577453527919715, 33.68082892595767, 35.22350436787768, 36.212613268842894, 38.08197656670742, 37.30408360112178, 37.95604884285448, 39.60721623670514, 40.264174065575624, 45.77534365433292, 57.25012682117401, 56.921762229040695, 52.83418534835231, 52.71217986093169, 53.140170990944604, 54.41220605747602, 56.49276287239014, 58.69780797961482, 60.897371283306335, 60.01163733629599, 62.32164248706019, 66.5080153471665, 77.64205104829045, 83.80644239037203, 93.6147531296434, 104.09680614062754, 99.14401453911385, 91.42833814682868, 89.87874155455575, 90.96141143308267, 94.15573561664038, 100.00369706373107, 108.06602180342581, 112.57476418518276, 114.9077981824693, 115.81341285585872, 120.60742590469337, 130.0096132082738, 141.08695909628977, 154.9758508976317, 169.2254112655649, 189.96423864768326, 205.79535472958864, 216.8617270913649, 225.7385757631245, 240.07582411195656, 248.11111797748617, 253.6691120390557, 257.7358354401678, 261.76377602027736, 262.9749545284158, 264.54363964321226, 264.46708081574485, 263.7219736663458, 262.9666561405128, 256.9916050968082, 253.36956899458457, 253.25480286956062, 253.35734687932916, 253.64214921830362, 253.66117111389616, 253.84242581929172, NaN, NaN, 23.96697483131655, 23.89003910957913, 24.477354445231256, 25.506191230228005, 26.901184895614865, 29.54876393697912, 31.384653743794107, 33.14558180129519, 34.68636869339689, 35.85889095256172, 36.66442014681849, 38.28040223046357, 41.21658371368227, 43.493428491811706, 45.991909824230426, 46.35541805476835, 43.631324268004484, 47.59572131620167, 55.607998971749176, 56.56654512641735, 50.42154817101768, 51.44467333287792, 58.05629929999922, 61.43483068953114, 62.974228234954936, 67.74977004169291, 65.90790158474151, 65.456956245275, 70.08316231408861, 77.13704248680268, 84.4047736668444, 89.75835036951288, 96.58526022683084, 102.38838933682752, 104.3009471879992, 102.26705422607986, 95.89027920968798, 95.59037538828518, 96.7003517105819, 97.42586875063795, 101.64162054528417, 109.8759487638304, 113.54403426794363, 117.38255388415831, 124.75385621421484, 138.01459628607387, 148.79660788660058, 159.7705768070378, 169.58448995411572, 180.24099126549658, 185.52871073344355, 199.18916884894327, 216.59993788489163, 233.77286885113293, 243.39179279006584, 247.05882278286467, 252.95068885117564, 256.21020245814964, 260.79848423572025, 262.84976695630974, 263.7068990183462, 263.36200705428564, 264.47666911381066, 260.38594550923847, 254.33263977190973, 252.53196777579336, 252.563463749937, 252.7395454627312, 252.90829948243402, 253.00336103489053, NaN, NaN, 21.195670453405842, 22.188916135029366, 23.84468442553567, 24.982391042121947, 26.08621539824771, 28.18082807625182, 29.243930291938494, 30.303790313269573, 31.143566906352177, 31.468935625804686, 32.89726479083633, 35.13542182624413, 37.115381996247535, 39.31703077430115, 41.81761420101114, 44.20281224264166, 46.99730677916215, 49.96946302093443, 51.9870405951668, 55.2596482209395, 55.36208942901638, 55.46401849150705, 60.41453325871219, 65.37141434995536, 61.95170812300536, 63.70954631779747, 63.70202712346572, 70.08734640163122, 72.84437483412111, 74.60728879080663, 81.65851432914495, 91.24039985812924, 97.62232222031535, 103.67878044041737, 109.19663028359317, 108.65982730615914, 113.1896717710949, 124.2245417525078, 126.56766350088466, 118.30581753648873, 123.31909364748486, 129.3658165421984, 134.5273628158968, 138.09117488120597, 145.7971191633128, 154.41286434922225, 168.69095213859794, 178.77205266829776, 196.62490287706288, 212.23765730759553, 227.9582624610713, 235.25937655620092, 239.5139578370475, 245.29373348512348, 249.44183520468562, 253.75132641167102, 256.7873980184183, 260.6507780103785, 261.7313348623411, 263.21850296252575, 264.0170144793085, 264.8415017786221, 264.6063162137331, 261.4610937242732, 253.97059248816254, 252.74138143019889, 253.06719810840985, 253.08621366281625, 253.28233864447057, NaN, NaN, 24.372857063040257, 24.370270771466448, 25.510779063415836, 26.280719230619937, 26.717963932115318, 27.967499951129707, 29.40057940757987, 31.681505668347555, 32.34289900608085, 34.291992817844246, 36.42653351390093, 38.29715581578848, 39.72668157276916, 42.04315249436061, 44.72656812848452, 47.25858769793706, 49.82988165785655, 52.36181768922954, 55.33108981986331, 59.109793823587864, 62.37292959399333, 63.47006330704947, 64.71290343406612, 66.98057955294188, 71.24018558438254, 74.32412844237798, 75.34670531876223, 72.4035660344671, 74.14975721474285, 75.68078948753491, 75.006689710218, 75.43666739083406, 78.88213121022946, 86.43556894654806, 93.33864312987546, 97.74245057890901, 95.6870925616293, 96.42152337905047, 103.98245416334774, 106.4886356356988, 106.87554642117236, 111.72726519645916, 119.54310237853859, 125.60646892608379, 127.55592930776105, 128.47265078117093, 135.588865493972, 143.86130592053925, 161.34492375945868, 174.26994523538778, 187.32686087168622, 198.08252238221925, 211.58201605490737, 225.40249765356623, 234.30238465880825, 241.34738963537995, 246.3832333376551, 252.03894626742203, 256.95891715961295, 261.49541718795825, 263.3507381790049, 263.1634448406584, 263.4037000126485, 261.99988175571747, 254.82818832662417, 252.1294389335514, 251.588101873147, 251.8327900437963, 252.07658316244923, 254.19743254436182, 255.25868899054007, 255.13073800330736, NaN, NaN, 253.7922838423942, 253.81747895562583, 253.84600804228634, 253.94078409694833, 253.94548179696878, 253.91521861049827, 253.923978697337, 254.01662736956325, 254.0840723573345, 252.91748258968482, 252.97496754136924, 253.40224075349477, 252.51708363892004, 252.579545295633, 252.45651352564414, 251.3347422480356, 251.565538102904, 216.6177812243208, 86.31386081935419, 61.58153836564415, 61.86084428637735, 65.74674464664233, 67.87087175894517, 69.33296964204763, 70.65639167776595, 73.88403641581742, 75.4848901247146, 77.2442953546329, 79.58584219048734, 82.88937080849597, 89.3353141230066, 94.76540462325362, 97.62564480952453, 99.39641974987522, 101.1576299358205, 104.0252502140031, 105.72447978051454, 105.89093163436402, 108.61953236752805, 113.10802345082419, 117.91919047976906, 128.03464775492657, 134.31978813936738, 141.3408495412661, 152.65231724041297, 169.4671256937398, 188.61437302860085, 200.7147427449083, 214.34154060052515, 224.6470242484939, 233.6891998403054, 242.7556271215318, 248.11908906401763, 251.48337881583595, 255.37795250414203, 259.4721820042675, 263.4726950631407, 264.4915238799946, 264.2257173362035, 256.24306423658044, 251.7958268711613, 251.36255878922748, 251.08657439801271, 250.76358529824083, 249.5340417664957, 249.1711959739924, 249.09940690996632, NaN, NaN, 24.922106606522696, 24.660119939866824, 24.72828509375323, 25.274414359102604, 25.709881377251087, 25.854047729663957, 26.88144011994814, 28.718020740999798, 29.116807030379434, 29.075104263751516, 30.097848198111826, 33.477765546969856, 37.00638967468955, 37.95784538359949, 38.42730649841856, 40.443371124691296, 44.33408760048329, 47.85819547096147, 50.67976876654289, 52.51220598737166, 52.063516288223596, 54.47962596895989, 60.4267706143667, 64.72501119910571, 67.3665723992014, 68.35238318106546, 69.22632788113887, 71.53694836756408, 73.52215750713286, 78.03288100225218, 79.35920262168139, 79.7903175553585, 80.33239277368149, 82.5319838393803, 85.836345010112, 88.80574928031058, 85.17578320681008, 83.19424927206282, 84.28600335222474, 96.28941424574691, 104.90548006776137, 110.37072277928185, 113.46606237276644, 124.21958190865891, 136.0221392910882, 143.26483442810496, 154.6496932559512, 165.78197555295068, 176.37253413166795, 185.49249073621934, 198.50651516669356, 214.6877017118266, 225.9509819433698, 236.01823343835272, 242.82772422762136, 248.9951445374831, 253.89641668828907, 256.5030070735777, 259.9323107720957, 263.3443531607177, 265.4930002322465, 265.50547890813004, 261.89182564580057, 252.96619544903388, 250.65531502328952, 250.84808391667227, 250.83042045731574, 250.0557267444252, 248.6783212604824, 248.64916094769035, NaN, NaN, 22.149384972008352, 22.296086300248813, 22.846643859023562, 23.872899380411447, 24.863950253501127, 27.625076447755667, 29.867948901625887, 31.18662168368748, 31.992568746594102, 33.49924938798738, 35.259901011594245, 37.16390049167275, 38.95718635015479, 39.20875388815881, 39.753858173035454, 44.01543368689123, 47.65990012473, 49.34762141308156, 51.287128178242114, 54.95450512247823, 58.03298564832189, 59.89799248829779, 62.20543246936147, 64.18871707667057, 65.29027932768835, 67.82965098521764, 71.58276603187147, 78.40922064454232, 82.70191918530826, 83.91623493262043, 85.90465439682771, 82.26011334819978, 84.00499129884301, 91.26540377987641, 94.79755085039213, 90.06234776608304, 90.7228131852584, 91.70549360873414, 98.42317796176263, 109.55054645173622, 113.86494117093417, 116.38047222177087, 116.84416813086527, 130.71675706778024, 143.26519364270086, 153.48914423643916, 168.93371055764408, 178.77672318881432, 188.31542897554567, 199.04359451357175, 211.47533977590396, 226.87858634168447, 238.25037363774624, 248.21892095925045, 251.492424069995, 255.79844566373376, 259.47439364590326, 262.29103776355873, 264.09397730784116, 266.0862273364447, 266.9851292441303, 260.58747860105984, 252.3501414578397, 251.57210156085318, 250.55045400478016, 249.86689594827055, 248.02442073311136, 246.48339395522353, 246.18053636838138, 246.5381472628425, NaN, NaN, 23.48784600631909, 23.5584175491109, 23.959601293150353, 25.022559918334288, 26.934282325414085, 29.285466896801577, 30.936933725148307, 32.44007136892288, 34.200617130727224, 35.81269254680137, 36.91013511797521, 36.978886140299366, 38.81114735609731, 41.014198547761445, 43.25217331838855, 45.5650194411642, 49.047287199177596, 50.547547322219884, 51.785253430912995, 55.196759459846106, 56.368063534964556, 58.49492122188108, 66.6424974676999, 70.76444934554063, 70.39797620584591, 70.83314643584458, 73.24559879696801, 77.71944261023148, 81.60630381762904, 81.9763078816847, 79.32932778792511, 77.64072842267787, 83.72280360377773, 86.36645937461056, 89.16058698284071, 93.34307951417581, 101.20746339373521, 103.65484191767139, 107.10105563106, 109.59304000093971, 113.37888715933346, 121.78682163711245, 134.22036354759447, 143.72640264482803, 154.26856435741067, 170.45811384056785, 187.29373436487546, 196.1866645749562, 214.27008078489675, 230.40566702417865, 241.55290895427817, 248.77300716655904, 254.28460721255857, 258.9195090674149, 263.7913146534133, 266.32097842658, 268.03655406201847, 267.418608037344, 261.8176500180895, 253.36929627738024, 250.59065186659652, 248.7244101304013, 247.6238900302599, 246.90316787520226, 246.51680291439493, 246.27171529430217, 245.97987825415808, NaN, NaN, 21.558805085169517, 21.482929647148413, 21.737933939148114, 22.507961183555707, 23.351388696272632, 25.668998901033216, 28.648776973191154, 31.62438710036343, 33.90256787329612, 34.89255133256194, 35.40288588098103, 36.610354901610144, 38.07536572476554, 39.02581873392504, 39.39165786069952, 40.45337433848972, 43.062812158070734, 47.03617445975762, 50.818320583978256, 53.901696500515804, 58.013573151548826, 61.462644287542965, 60.206491072494636, 58.28997140741683, 62.32896967144364, 69.599613216701, 71.21774805493676, 72.31966469618224, 74.59254827307798, 76.19584503976508, 79.86135507233533, 85.31211771189999, 84.51936151302277, 81.57560436940285, 83.62402800318672, 85.67001849277949, 89.48126489954919, 88.58670432275588, 90.48295323849099, 98.49000243756578, 100.0071081358469, 105.52977078073691, 113.44020517692184, 117.86184348832136, 128.93202853023092, 138.73261678657593, 147.7719794944494, 154.9862613879334, 160.05278279525496, 168.61273745171187, 178.28970939151267, 192.99710725271012, 204.7149850624625, 224.8423675195162, 238.77300944300157, 245.50840437219702, 249.85554637457753, 254.49000845869566, 258.6723480008297, 262.1512689948434, 266.88506085235605, 267.77543434063836, 261.0617280290614, 253.74935329681102, 249.49062894198843, 248.96871635361305, 249.44206946090347, 249.34853363169134, 248.84052178609983, 247.60465903358946, 247.17184282107067, NaN, NaN, 21.303711350666205, 21.33775956932482, 21.887092633765374, 23.35694355873693, 24.824756615240325, 27.43243991944322, 30.37420620200196, 31.839554384243275, 33.30872285639525, 34.63214538622534, 35.548809700198746, 36.390663325533424, 37.081844115758415, 38.105087996601995, 40.162890874888454, 41.5557524057735, 42.06741072023655, 43.46111753802166, 45.294303964432, 47.97228042803912, 50.17668635584313, 53.18293591966205, 58.61043683730525, 63.00780359521036, 64.7652426682247, 68.0667089993597, 65.79403743359683, 69.08814469850753, 71.95217385030493, 73.3468914960999, 74.29984466599531, 77.38211087076412, 80.31008980589759, 85.07796061207537, 90.3635639776416, 91.98580559050536, 87.42739692863508, 87.19894797468709, 91.52811055029838, 95.56746839132263, 96.14972247960293, 104.51511929519108, 108.47973432556661, 111.12585729142769, 115.09528346789656, 118.07707764687504, 122.17878363627192, 124.22403667918528, 131.6543302922779, 144.84124635564942, 150.86315939868166, 163.8855688691145, 177.49551586080972, 189.1039348788173, 199.71632524657204, 205.2815277002312, 211.7936054408003, 219.82810280305907, 230.1034953511598, 238.80800030230247, 243.8177793121005, 248.88526495352545, 254.8785681538595, 260.6527807948851, 262.66400896538113, 262.5356959556318, 259.9411316688745, 251.81985915441928, 249.10166821696367, 249.34696404561026, 249.60279491475262, 249.64278545995109, 249.09367928911777, NaN, NaN, 22.924291215877044, 22.2954986257626, 22.623017891066453, 25.56416756665099, 29.499803815722803, 32.072677786245535, 32.98714042427955, 32.8339445731035, 33.49259818970274, 33.891024304951685, 35.98367129014639, 37.96277590894452, 39.428876347090636, 41.81398203531724, 43.13458598022031, 44.45411327039092, 46.47099406064557, 48.41399282369985, 52.59786903094238, 55.56915830144296, 59.381962854933, 65.32918405619307, 68.96118243800049, 70.38656515331851, 69.167598907388, 67.61926464338575, 73.33928680760398, 78.19409549875898, 81.9442048031078, 83.92580327289825, 84.35315632960388, 86.32754635006883, 92.50673018128607, 93.05537238449057, 94.48634781824907, 94.93283490351148, 99.55142033238361, 100.20291448481429, 96.24353915938228, 107.71068157347537, 117.31765517069717, 122.05234873296021, 121.93589761519324, 127.85825789175274, 141.75417135800035, 150.3958333633047, 164.44420916170958, 175.1412619040059, 183.9001240043914, 193.59607302887963, 202.55782698410997, 213.49684744397746, 222.22757681863865, 231.43810624186048, 240.71042231349483, 245.99125290527547, 248.9851683971997, 251.7952363503293, 258.24085648605796, 261.1303789882261, 262.82192198847315, 263.94003487192805, 262.4767115575069, 252.47229985449658, 249.58936549096703, 249.44369372734042, 249.41020622144887, 249.05827868092518, 248.11553719810274, 247.89491858395857, NaN, NaN, 25.652841532401624, 25.206326012576746, 26.455131705447098, 28.36563643502997, 29.98246568910988, 31.15508896483024, 32.03253223120575, 33.09293798691342, 34.15643495956283, 35.36405124884207, 35.94636317840649, 35.94104421435955, 37.51588376770436, 39.420770249279514, 41.327169937942706, 43.26994786958847, 43.592225064792345, 44.17443953574209, 46.78206542660271, 49.45625366349167, 51.40176799606656, 53.30657372876148, 57.85056131416775, 64.38320308549328, 69.44200659062275, 73.47564570759249, 71.63853276715965, 71.56429855499582, 75.31618059647151, 83.01924637988897, 87.6429946308429, 88.75644985046935, 90.67070122900316, 93.30305511595235, 95.28891969266365, 96.98112961951922, 99.19138603577906, 100.22917039334077, 105.00885826047742, 110.89772849685595, 110.21941677827024, 122.52655100526617, 142.97930457744368, 151.92232663947408, 162.29253548018534, 175.71045083797654, 191.52280495832497, 205.90669099007525, 216.57797432574304, 229.03136084538193, 239.44029780517556, 245.54633375945, 249.91466538453872, 254.9929271562293, 262.2867121601881, 265.57616353045364, 264.56496807696107, 263.3008172165738, 261.6562560699711, 260.10092550766234, 256.2453106408829, 254.03231485209483, 252.0599256726362, 249.3484359787459, 248.07596120426058, 248.18718068457403, 248.41912149891667, NaN, NaN, 24.39443915664378, 23.83793795939749, 24.75645701910413, 26.48292507683478, 28.2096449431594, 29.863224908564554, 32.21627997061758, 33.24491383418324, 33.828249775735344, 35.07498487835386, 35.328720362076055, 36.27844062308614, 38.47769068913537, 40.05193013607993, 42.031754141963695, 43.45480206300818, 43.37215004560782, 44.172380976896925, 45.45002544193958, 47.79487772015818, 50.87592767791967, 53.51638618130603, 56.07734524481222, 59.22895560623408, 64.94863929503592, 69.12876938315902, 72.1369039522421, 70.3002047444545, 66.10708402704192, 68.5292396335672, 71.17004575743836, 74.68217423966868, 81.20323015509595, 85.53251294985971, 87.14424558591163, 90.52877755055128, 93.39004892223606, 94.27558922971645, 96.61956983502064, 99.27451196225049, 102.1531360994222, 106.02841306359558, 108.98688500788533, 116.00311175558905, 137.16000781997298, 151.606919738498, 164.67141702847445, 186.82262576168378, 203.61589651286877, 213.0546257457534, 219.82550987947567, 228.08888115627119, 237.32410750859034, 243.79613579509896, 249.0950087539343, 253.32986808960212, 258.3844841424484, 262.6070564335954, 264.06769870237844, 263.6732272553881, 262.69192417664215, 260.840985037835, 257.3022323512535, 252.84926774487462, 250.91450794971507, 250.37970114274964, 250.24922832690802, 250.42868382812628, NaN, NaN, 25.870775190580165, 25.61027627552401, 26.084526543163136, 26.41065761282741, 26.184499193271705, 27.909794398975183, 28.898186818908695, 31.43542044255447, 32.39156476449624, 33.08542355557211, 34.589695581581374, 36.75629407499566, 38.958092779202865, 41.34240903338128, 43.21309280706205, 44.60776862585186, 46.03561123836557, 47.830303462714795, 50.57991235712032, 52.70351204812094, 53.50050339299118, 55.25231916612455, 59.06267361264662, 64.56068050241304, 69.10854667389148, 71.83299226457656, 69.91194816249664, 69.75375129886274, 69.89347254819715, 70.4792393776912, 75.0193947726804, 77.58353979580754, 83.74665660550767, 87.0492963138433, 90.13720287445227, 95.64901345083065, 96.89750527046135, 99.85771125076072, 97.75056807698688, 98.33507227700994, 105.42804340773995, 107.21356224056031, 118.69443386899866, 135.7767605200206, 150.6964459431458, 157.0875406097836, 165.91229761442438, 183.48233728161884, 199.12013017034164, 210.08996794314152, 219.29315493965737, 228.44852786502568, 235.1868933990256, 239.03360589678607, 245.45714922704204, 250.4671419917587, 255.30376062275582, 258.03282461228974, 260.3885082288746, 263.6998922598336, 264.3651716012192, 265.1578302888916, 264.6641952673486, 261.7055063163389, 256.3466794653368, 253.21326076837627, 250.52082587832092, 249.91749939502452, 249.82973892722484, NaN, NaN, 24.06048202797541, 21.62606452724144, 20.59097679389164, 21.323826746638336, 22.71940207456684, 23.96646477352765, 25.656537241745156, 26.314935727339098, 27.563208235240516, 28.956875790774287, 30.8645434051679, 32.846866348545014, 33.652560196814434, 35.0474221733259, 37.39774621951811, 42.09848798311983, 43.786547597146104, 45.400923048383646, 47.52855404006613, 50.82844523728666, 51.92440464204934, 53.685052002946456, 55.953045933678574, 63.953735602762954, 68.50930038957291, 71.23346759230179, 72.39723357676633, 71.44000364556778, 70.55514654800504, 70.77128262258128, 75.61478530563907, 81.1929136359639, 84.4200411576779, 89.0372812265571, 91.07832379764324, 93.50062669238886, 95.25212712492696, 98.64097326960899, 100.56039855197058, 100.11897163653256, 101.29847004085859, 94.9959139669918, 98.5030688809473, 106.73063499661889, 110.39690111276609, 124.41586936409105, 140.19782997557505, 155.44683220996805, 164.95729010535544, 175.25894688975924, 190.88058464006346, 204.16596099620222, 210.96298875520975, 220.56796005275825, 229.88538292764017, 236.18655886795418, 239.24559382536393, 246.09827742870002, 251.10763141649045, 254.25880313136406, 255.8940261993349, 260.0221358817254, 262.81802655436144, 264.48117472407864, 265.0549914257371, 264.5506749763318, 263.49583654650553, 255.88761243159743, 250.58070711663473, 249.82190071102448, 250.1366970659754, 250.25103172917932, NaN, NaN, 19.157434829515488, 19.007121432430697, 20.698682968966345, 21.72584862234667, 21.571180700901262, 22.15426928604878, 23.916889297863843, 25.975514198683758, 27.592059309337245, 28.542780822956516, 30.374897749768156, 32.064042743722176, 33.23717997598079, 37.57164721990669, 42.56709016161002, 45.067246065551174, 47.12144606815711, 47.928536025203414, 50.78556126551974, 54.89520996945702, 56.98292968938007, 61.38257430165334, 65.19770035086616, 67.83110564033787, 71.20659911218104, 72.80899344064717, 73.75772520605578, 76.03149997870757, 73.53634581849289, 78.81665276762175, 86.74222108683095, 90.85332661983028, 93.26624711254607, 95.69331937604113, 101.29546344029826, 104.6739537688777, 103.21290070147822, 101.31454584921964, 99.70551530696302, 108.82303824248109, 114.64006514741794, 117.29434537814149, 126.74825916453965, 136.92695285616588, 153.024432150888, 164.27757287768554, 171.89011545049695, 184.55721982511972, 197.7627792351771, 209.44714879883742, 223.9336666342261, 232.0223913200024, 240.17178778648056, 245.4002055995207, 247.37086480876206, 248.45778234048356, 253.6207805860712, 256.8013399397391, 259.7238663485176, 262.1241001975999, 262.6571937095781, 262.91446116634626, 262.54382050287273, 258.8954159027256, 252.89231824797633, 250.34764423646857, 249.74444061228482, 249.91827787317658, 250.02169653834437, 250.14190206234107, NaN, NaN, 19.560556519126795, 19.18971312907147, 19.73848255684189, 21.206902482706163, 21.573128332582503, 22.267302234453005, 23.32978797076494, 24.57596392634873, 25.491092581126406, 26.000311335011858, 27.134783557717494, 29.411855478183348, 30.91793442466482, 33.156690990500785, 36.425743695456525, 38.36798609296721, 40.67912094958336, 43.0667165761046, 45.81763563493848, 48.018469356808666, 49.89161154064356, 51.43384283317056, 57.04613676403616, 63.543750274626795, 67.3921357480692, 71.13139665577246, 72.56427542033748, 75.53206360937959, 78.38730653332964, 80.46974009053919, 83.88281239328093, 85.96907739163952, 94.88836211322862, 102.59422255019098, 107.86852350230504, 112.70451897770343, 124.70287960172449, 128.66046734340043, 130.1898596810392, 132.82491892339286, 119.00546473332706, 109.92204522165245, 121.68834586126651, 127.76058162857144, 137.79326821189332, 143.256430219739, 154.787399203126, 163.9880877673297, 174.18242483028905, 190.67090820944696, 204.59292388951954, 212.53338886633193, 218.96729195929655, 234.04857734336437, 244.6049571142893, 247.19847968318444, 254.38270004668988, 257.8788289457661, 261.18422327216655, 262.83969054222354, 264.01199737796964, 263.27741378169753, 256.1053884596102, 251.53924893711692, 250.49194632655153, 250.53193319301946, 250.35424730794517, 250.2572081628754, 250.67477787968866, 250.80111928496865, NaN, NaN, 22.624691872554713, 22.3643122996152, 22.546783285814122, 23.021764246479954, 22.870216530897423, 25.847295743174275, 27.428502238878156, 28.78388949293049, 29.992755070201703, 30.867980450815345, 32.51588159948183, 34.535156467643844, 36.11115348068115, 37.94294319921429, 39.587134985067664, 41.01042434967362, 42.764180622829784, 44.337897737914446, 45.363485286700886, 46.569707047354775, 48.692873608095766, 51.259530439566355, 55.47300319895375, 60.05508811559973, 65.37362267413434, 68.30850930345642, 70.69200691369939, 72.52413829933879, 77.28815890671991, 81.13548382040183, 84.07395601517413, 84.80306148176354, 87.73101771729277, 92.85839329067332, 105.33202391852318, 125.70200962114743, 127.72549428600657, 132.871578963824, 138.21045277257303, 138.79253373519398, 143.2050043748133, 146.91750451963017, 148.4465097909897, 160.49339956460187, 167.2907687433464, 182.63691510690853, 200.369188670614, 208.43725975328272, 212.62259150439976, 218.1021840964203, 224.7338832418125, 236.36462176321874, 244.23099815342366, 248.83282897494786, 252.92458437775358, 257.78955230350033, 260.20385631574055, 262.62120770817046, 265.90735969682925, 262.8183666647025, 256.6403519752979, 252.62887803005802, 252.18597563612119, 252.51791436046338, 252.28151763719382, 250.99268165479413, 250.2744650727306, 250.17185083862626, NaN}
    PARAMETERS =   "CHLA",   "DENSITY",   "DOXY"
    DOXY_QC = 
      {9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9, 9, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 9}
    CHLA_INSTRUMENT = 
      {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
    DOXY_INSTRUMENT = 
      {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
}

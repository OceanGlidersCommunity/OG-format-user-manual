netcdf file:/Users/sevadjian/projects/sushi/missions_netcdf/mission_output/OG-10-202400415/20240607/sp028_20230202T1637_R.nc {
  dimensions:
    n_measurements = UNLIMITED;   // (372 currently)
  variables:
    String trajectory;
      :cf_role = "trajectory_id";
      :comment = "A trajectory is one deployment of a glider. The format is platform_id-YYYYMMDDThhmm. Where the time is the start of the first dive of the trajectory.";
      :long_name = "Trajectory Name";

    int profile_index(n_measurements=372);
      :comment = "Sequential profile number within the trajectory, extended for use along the n_measurements dimension. Use this variable for indexing or shaping the data. The first profile has a value of 1 and is incremented for each successive profile contained in the trajectory.";
      :ioos_category = "Identifier";
      :long_name = "Profile Number";
      :valid_max = 2147483647; // int
      :valid_min = 1; // int
      :_FillValue = -999; // int
      :_ChunkSizes = 1024U; // uint

    double time_profile(n_measurements=372);
      :_CoordinateAxisType = "Time";
      :long_name = "Profile Time";
      :axis = "T";
      :calendar = "gregorian";
      :comment = "An estimate of the time of the mid-point of each profile. time_profile = time_gps + 0.75 * (time_gps_end - time_gps);";
      :ioos_category = "Time";
      :observation_type = "calculated";
      :platform = "platform_meta";
      :standard_name = "time";
      :time_origin = "01-JAN-1970 00:00:00";
      :units = "seconds since 1970-01-01T00:00:00Z";
      :ancillary_variables = "time_profile_qc";
      :_ChunkSizes = 512U; // uint

    int time_profile_qc(n_measurements=372);
      :_FillValue = -127; // int
      :long_name = "Profile Time Quality Flag";
      :standard_name = "aggregate_quality_flag";
      :valid_max = 9; // int
      :valid_min = 0; // int
      :flag_values = 1, 2, 3, 4, 9; // int
      :flag_meanings = "good not_evaluated questionable bad missing";
      :comment = "1=Good/Pass, 2=Not Evaluated, 3=Questionable, Suspect or of High Interest, 4=Fail/Bad, 9=Missing Data. See the references for more details on the flag meanings.";
      :references = "Paris. Intergovernmental Oceanographic Commission of UNESCO, 2013. Ocean Data Standards, Vol.3:Recommendation for a Quality Flag Scheme for the Exchange of Oceanographic and Marine    Meteorological Data. (IOC Manuals and Guides, 54, Vol. 3.) 12 pp. (English.)(IOC/2013/MG/54-3) https://repository.oceanbestpractices.org/bitstream/handle/11329/413/MG54_3.doc";
      :_ChunkSizes = 372U; // uint

    double latitude_profile(n_measurements=372);
      :_FillValue = -999.0; // double
      :_CoordinateAxisType = "Lat";
      :long_name = "Profile Latitude, Mid-Point";
      :axis = "Y";
      :colorBarMaximum = 90.0; // double
      :colorBarMinimum = -90.0; // double
      :comment = "An estimate of the latitude at the mid-point of each profile. latitude_profile = latitude_gps + 0.75 * (latitude_gps_end - latitude_gps);";
      :ioos_category = "Location";
      :observation_type = "calculated";
      :platform = "platform_meta";
      :standard_name = "latitude";
      :units = "degrees_north";
      :valid_max = 90.0; // double
      :valid_min = -90.0; // double
      :ancillary_variables = "latitude_profile_qc";
      :_ChunkSizes = 372U; // uint

    int latitude_profile_qc(n_measurements=372);
      :_FillValue = -127; // int
      :long_name = "Profile Latitude Mid-Point Quality Flag";
      :standard_name = "aggregate_quality_flag";
      :valid_max = 9; // int
      :valid_min = 0; // int
      :flag_values = 1, 2, 3, 4, 9; // int
      :flag_meanings = "good not_evaluated questionable bad missing";
      :comment = "1=Good/Pass, 2=Not Evaluated, 3=Questionable, Suspect or of High Interest, 4=Fail/Bad, 9=Missing Data. See the references for more details on the flag meanings.";
      :references = "Paris. Intergovernmental Oceanographic Commission of UNESCO, 2013. Ocean Data Standards, Vol.3:Recommendation for a Quality Flag Scheme for the Exchange of Oceanographic and Marine    Meteorological Data. (IOC Manuals and Guides, 54, Vol. 3.) 12 pp. (English.)(IOC/2013/MG/54-3) https://repository.oceanbestpractices.org/bitstream/handle/11329/413/MG54_3.doc";
      :_ChunkSizes = 372U; // uint

    double latitude_uv(n_measurements=372);
      :_FillValue = -999.0; // double
      :long_name = "Latitude of Underwater Segment Mid-Point Estimate";
      :axis = "Y";
      :colorBarMaximum = 90.0; // double
      :colorBarMinimum = -90.0; // double
      :comment = "This latitude variable is provided specifically for use with the depth-averaged current variables u and v. The value is an estimate of the glider location at the midpoint of the underwater segment. It differs from the latitude variable which is the estimate of the mid-point of the profile which is at 3/4 of the underwater segment. The value is interpolated to provide an estimate of the mid-point of the entire underwater segment, which may consist of 1 or more dives. Calculated using surface GPS positions at the start and end of the dive. Where, latitude_uv = latitude_gps + 0.5 * (latitude_gps_end - latitude_gps);";
      :ioos_category = "Location";
      :observation_type = "calculated";
      :platform = "platform_meta";
      :standard_name = "latitude";
      :units = "degrees_north";
      :valid_max = 90.0; // double
      :valid_min = -90.0; // double
      :ancillary_variables = "latitude_uv_qc";
      :_ChunkSizes = 372U; // uint

    int latitude_uv_qc(n_measurements=372);
      :_FillValue = -127; // int
      :long_name = "Latitude of Underwater Segment Mid-Point Estimate Quality Flag";
      :valid_max = 9; // int
      :valid_min = 1; // int
      :flag_values = 1, 2, 3, 4, 9; // int
      :flag_meanings = "good not_evaluated questionable bad missing";
      :comment = "1=Good/Pass, 2=Not Evaluated, 3=Questionable, Suspect or of High Interest, 4=Fail/Bad, 9=Missing Data. See the references for more details on the flag meanings.";
      :references = "Paris. Intergovernmental Oceanographic Commission of UNESCO, 2013. Ocean Data Standards, Vol.3:Recommendation for a Quality Flag Scheme for the Exchange of Oceanographic and Marine    Meteorological Data. (IOC Manuals and Guides, 54, Vol. 3.) 12 pp. (English.)(IOC/2013/MG/54-3) https://repository.oceanbestpractices.org/bitstream/handle/11329/413/MG54_3.doc";
      :_ChunkSizes = 372U; // uint

    double longitude_profile(n_measurements=372);
      :_FillValue = -999.0; // double
      :long_name = "Profile Mid-Point Longitude";
      :axis = "X";
      :comment = "An estimate of the longitude at the mid-point of each profile. longitude_profile = longitude_gps + 0.75 * (longitude_gps_end - longitude_gps);";
      :ioos_category = "Location";
      :observation_type = "calculated";
      :platform = "platform_meta";
      :standard_name = "longitude";
      :units = "degrees_east";
      :valid_max = 180.0; // double
      :valid_min = -180.0; // double
      :ancillary_variables = "longitude_profile_qc";
      :_ChunkSizes = 372U; // uint

    int longitude_profile_qc(n_measurements=372);
      :_FillValue = -127; // int
      :long_name = "Profile Longitude Quality Flag";
      :standard_name = "aggregate_quality_flag";
      :valid_max = 9; // int
      :valid_min = 1; // int
      :flag_values = 1, 2, 3, 4, 9; // int
      :flag_meanings = "good not_evaluated questionable bad missing";
      :comment = "1=Good/Pass, 2=Not Evaluated, 3=Questionable, Suspect or of High Interest, 4=Fail/Bad, 9=Missing Data. See the references for more details on the flag meanings.";
      :references = "Paris. Intergovernmental Oceanographic Commission of UNESCO, 2013. Ocean Data Standards, Vol.3:Recommendation for a Quality Flag Scheme for the Exchange of Oceanographic and Marine    Meteorological Data. (IOC Manuals and Guides, 54, Vol. 3.) 12 pp. (English.)(IOC/2013/MG/54-3) https://repository.oceanbestpractices.org/bitstream/handle/11329/413/MG54_3.doc";
      :_ChunkSizes = 372U; // uint

    double longitude_uv(n_measurements=372);
      :_FillValue = -999.0; // double
      :long_name = "Longitude of Underwater Segment (Mid-Point Estimate)";
      :axis = "X";
      :comment = "This longitude variable is provided specifically for use with the depth-averaged current variables u and v. The value is an estimate of the glider location at the midpoint of the underwater segment. It differs from the longitude_profile variable which is the estimate of the mid-point of the profile which is at 3/4 of the underwater segment. The value is interpolated to provide an estimate of the mid-point of the entire underwater segment, which may consist of 1 or more dives. Calculated using surface GPS positions at the starta nd end of the dive. Where, longitude_uv = longitude_gps + 0.5 * (longitude_gps_end - longitude_gps);";
      :ioos_category = "Location";
      :observation_type = "calculated";
      :platform = "platform_meta";
      :standard_name = "longitude";
      :units = "degrees_east";
      :valid_max = 180.0; // double
      :valid_min = -180.0; // double
      :ancillary_variables = "longitude_uv_qc";
      :_ChunkSizes = 372U; // uint

    int longitude_uv_qc(n_measurements=372);
      :_FillValue = -127; // int
      :long_name = "Longitude of Underwater Segment (Mid-Point Estimate) Quality Flag";
      :valid_max = 9; // int
      :valid_min = 1; // int
      :flag_values = 1, 2, 3, 4, 9; // int
      :flag_meanings = "good not_evaluated questionable bad missing";
      :comment = "1=Good/Pass, 2=Not Evaluated, 3=Questionable, Suspect or of High Interest, 4=Fail/Bad, 9=Missing Data. See the references for more details on the flag meanings.";
      :references = "Paris. Intergovernmental Oceanographic Commission of UNESCO, 2013. Ocean Data Standards, Vol.3:Recommendation for a Quality Flag Scheme for the Exchange of Oceanographic and Marine    Meteorological Data. (IOC Manuals and Guides, 54, Vol. 3.) 12 pp. (English.)(IOC/2013/MG/54-3) https://repository.oceanbestpractices.org/bitstream/handle/11329/413/MG54_3.doc";
      :_ChunkSizes = 372U; // uint

    double time_uv(n_measurements=372);
      :_FillValue = -999.0; // double
      :long_name = "Time Estimate for Underwater Segment";
      :axis = "T";
      :comment = "This time variable is provided for use with the depth-averaged current variables u and v. The value is an estimate of the glider location at the midpoint of the underwater segment. The value is interpolated to provide an estimate of the mid-point of the entire underwater segment, which may consist of 1 or more dives. Calculated using surface GPS times at the start and end of the dive. Where, time_uv = time_gps + 0.5 * (time_gps_end - time_gps);";
      :ioos_category = "Time";
      :observation_type = "calculated";
      :platform = "platform_meta";
      :standard_name = "time";
      :units = "seconds since 1970-01-01T00:00:00Z";
      :time_origin = "01-JAN-1970 00:00:00";
      :ancillary_variables = "time_uv_qc";
      :_ChunkSizes = 372U; // uint

    int time_uv_qc(n_measurements=372);
      :_FillValue = -127; // int
      :coverage_content_type = "qualityInformation";
      :long_name = "Time Estimate for Underwater Segment Quality Flag";
      :valid_max = 9; // int
      :valid_min = 1; // int
      :flag_values = 1, 2, 3, 4, 9; // int
      :flag_meanings = "good not_evaluated questionable bad missing";
      :comment = "1=Good/Pass, 2=Not Evaluated, 3=Questionable, Suspect or of High Interest, 4=Fail/Bad, 9=Missing Data. See the references for more details on the flag meanings.";
      :references = "Paris. Intergovernmental Oceanographic Commission of UNESCO, 2013. Ocean Data Standards, Vol.3:Recommendation for a Quality Flag Scheme for the Exchange of Oceanographic and Marine    Meteorological Data. (IOC Manuals and Guides, 54, Vol. 3.) 12 pp. (English.)(IOC/2013/MG/54-3) https://repository.oceanbestpractices.org/bitstream/handle/11329/413/MG54_3.doc";
      :_ChunkSizes = 372U; // uint

    double time(n_measurements=372);
      :_FillValue = -999.0; // double
      :_CoordinateAxisType = "Time";
      :long_name = "Time of Each Observation";
      :axis = "T";
      :calendar = "gregorian";
      :comment = "Time stamp at each point in the underwater profile during a dive. This time stamp corresponds to the acquisition of the sensor data.";
      :ioos_category = "Time";
      :observation_type = "measured";
      :platform = "platform_meta";
      :standard_name = "time";
      :time_origin = "01-JAN-1970 00:00:00";
      :units = "seconds since 1970-01-01T00:00:00Z";
      :_ChunkSizes = 372U; // uint

    int time_qc(n_measurements=372);
      :_FillValue = -127; // int
      :comment = "Subsurface time values are more accurate than subsurface latitude and longitude. Subsurface positions are best estimates with lower accuracy. See the corresponding position variable metadata for more details. 1=Good/Pass, 2=Not Evaluated, 3=Questionable, Suspect or of High Interest, 4=Fail/Bad, 9=Missing Data. See the references for more details on the flag meanings.";
      :coverage_content_type = "qualityInformation";
      :flag_values = 1, 2, 3, 4, 9; // int
      :flag_meanings = "good not_evaluated questionable bad missing";
      :long_name = "Quality Flag for the Time of Each Observation";
      :standard_name = "aggregate_quality_flag";
      :references = "Paris. Intergovernmental Oceanographic Commission of UNESCO, 2013. Ocean Data Standards, Vol.3:Recommendation for a Quality Flag Scheme for the Exchange of Oceanographic and Marine    Meteorological Data. (IOC Manuals and Guides, 54, Vol. 3.) 12 pp. (English.)(IOC/2013/MG/54-3) https://repository.oceanbestpractices.org/bitstream/handle/11329/413/MG54_3.doc";
      :valid_max = 9; // int
      :valid_min = 0; // int
      :_ChunkSizes = 372U; // uint

    double wcur_x(n_measurements=372);
      :_FillValue = -999.0; // double
      :ancillary_variables = "wcur_qc wcur_qc_tests";
      :colorBarMaximum = 0.5; // double
      :colorBarMinimum = 0.5; // double
      :comment = "The depth-averaged current is an estimate of the net current measured while the glider is underwater. The value is calculated over the entire underwater segment. The latitude_uv, longitude_uv and time_uv variables provide the location and time for this variable. Additional velocity data are available from the acoustic doppler current profiler (ADCP). Please contact us at idgdata@ucsd.edu if you are interested in the ADCP data.";
      :coordinates = "time_uv longitude_uv latitude_uv";
      :coverage_content_type = "physicalMeasurement";
      :ioos_category = "Location";
      :long_name = "U, Depth-Averaged Eastward Sea Water Velocity";
      :observation_type = "calculated";
      :platform = "platform_meta";
      :standard_name = "eastward_sea_water_velocity";
      :units = "m s-1";
      :valid_max = 10.0; // double
      :valid_min = -10.0; // double
      :vocabulary = "https://vocab.nerc.ac.uk/collection/OG1/current";
      :_ChunkSizes = 372U; // uint

    double wcur_y(n_measurements=372);
      :_FillValue = -999.0; // double
      :ancillary_variables = "wcur_qc wcur_qc_tests";
      :colorBarMaximum = 0.5; // double
      :colorBarMinimum = 0.5; // double
      :comment = "The depth-averaged current is an estimate of the net current measured while the glider is underwater. The value is calculated over the entire underwater segment. The latitude_uv, longitude_uv and time_uv variables provide the location and time for this variable. Additional velocity data are available from the acoustic doppler current profiler (ADCP). Please contact us at idgdata@ucsd.edu if you are interested in the ADCP data.";
      :coordinates = "time_uv longitude_uv latitude_uv";
      :coverage_content_type = "physicalMeasurement";
      :ioos_category = "Location";
      :long_name = "V, Depth-Averaged Northward Sea Water Velocity";
      :observation_type = "calculated";
      :platform = "platform_meta";
      :standard_name = "northward_sea_water_velocity";
      :units = "m s-1";
      :valid_max = 10.0; // double
      :valid_min = -10.0; // double
      :vocabulary = "https://vocab.nerc.ac.uk/collection/OG1/current";
      :_ChunkSizes = 372U; // uint

    int wcur_qc(n_measurements=372);
      :_FillValue = -127; // int
      :comment = "The depth averaged velocity calculation is dependent on the glider position at the start and end of each dive. These flags are derived from the GPS flags for the dive. 1=Good/Pass, 2=Not Evaluated, 3=Questionable, Suspect or of High Interest, 4=Fail/Bad, 9=Missing Data. See the references for more details on the flag meanings.";
      :coverage_content_type = "qualityInformation";
      :flag_values = 1, 2, 3, 4, 9; // int
      :flag_meanings = "good not_evaluated questionable bad missing";
      :long_name = "Depth-Averaged Sea Water Velocity Quality Flag";
      :standard_name = "aggregate_quality_flag";
      :valid_max = 9; // int
      :valid_min = 1; // int
      :_ChunkSizes = 372U; // uint

    int wcur_qc_tests(n_measurements=372);
      :_FillValue = -127; // int
      :coverage_content_type = "qualityInformation";
      :long_name = "Depth-Averaged Eastward Sea Water Velocity Quality Flag";
      :valid_max = 99; // int
      :valid_min = 0; // int
      :flag_values = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 99; // int
      :flag_meanings = "gps_good gps_day_problem gps_repeat gps_backward gps_too_fast_on_surface gps_too_soon gps_too_far gps_bad_hdop gps_bad_status gps_no_surfacing gps_manual gps_no_dive";
      :standard_name = "quality_flag";
      :comment = "The depth averaged velocity calculation on the glider position at the start and end of each dive. These flags are derived from the GPS flags for the dive. gps_good=0 gps_day_problem=1 gps_repeat=2 gps_backward=3 gps_too_fast_on_surface=4 gps_too_soon=5 gps_too_far=6 gps_bad_hdop=7 gps_bad_status=8 gps_no_surfacing=9 gps_manual=10 gps_no_dive=99";
      :_ChunkSizes = 372U; // uint

    double depth(n_measurements=372);
      :_FillValue = -999.0; // double
      :_CoordinateAxisType = "Height";
      :_CoordinateZisPositive = "down";
      :ancillary_variables = "depth_qc";
      :axis = "Z";
      :colorBarMaximum = 2000.0; // double
      :colorBarMinimum = 0.0; // double
      :colorBarPalette = "OceanDepth";
      :ioos_category = "Location";
      :long_name = "Depth";
      :observation_type = "calculated";
      :platform = "platform_meta";
      :positive = "down";
      :reference_datum = "sea-surface";
      :sensor = "sensor_ctd";
      :standard_name = "depth";
      :units = "m";
      :valid_max = 2000.0; // double
      :valid_min = 0.0; // double
      :vocabulary = "https://vocab.nerc.ac.uk/collection/OG1/current";
      :comment = "Depth values are calculated from pressure. A Spray glider profiles on the ascent, collecting sensor data beginning in deeper water and ending at the surface.";
      :_ChunkSizes = 372U; // uint

    int depth_qc(n_measurements=372);
      :_FillValue = -127; // int
      :comment = "1=Good/Pass, 2=Not Evaluated, 3=Questionable, Suspect or of High Interest, 4=Fail/Bad, 9=Missing Data. See the references for more details on the flag meanings.";
      :coverage_content_type = "qualityInformation";
      :long_name = "Depth Quality Flag";
      :standard_name = "aggregate_quality_flag";
      :flag_values = 1, 2, 3, 4, 9; // int
      :flag_meanings = "good not_evaluated questionable bad missing";
      :references = "Paris. Intergovernmental Oceanographic Commission of UNESCO, 2013. Ocean Data Standards, Vol.3:Recommendation for a Quality Flag Scheme for the Exchange of Oceanographic and Marine    Meteorological Data. (IOC Manuals and Guides, 54, Vol. 3.) 12 pp. (English.)(IOC/2013/MG/54-3) https://repository.oceanbestpractices.org/bitstream/handle/11329/413/MG54_3.doc";
      :valid_max = 9; // int
      :valid_min = 0; // int
      :_ChunkSizes = 372U; // uint

    double latitude(n_measurements=372);
      :_FillValue = -999.0; // double
      :long_name = "Estimated Subsurface Latitude";
      :colorBarMaximum = 90.0; // double
      :colorBarMinimum = -90.0; // double
      :comment = "Estimated position of the glider underwater during a dive. Use the GPS position variables for accurate positions at the surface. Use caution with these estimated subsurface position values, the deviation from actual position may be several hundreds of meters! Estimations are a dead reckoning using the GPS positions at the start and end of the dive, and the gliders estimated velocity. The calculation methods are described in: \'Rudnick, D. L., Sherman, J. T., & Wu, A. P. (2018). Depth-average velocity from Spray underwater gliders. Journal of Atmospheric and Oceanic Technology, (2018), 35, 1665-1673; doi: https://doi.org/10.1175/JTECH-D-17-0200.1\'. The accuracy attribute reflects an accuracy of approximately +/-800m (0.007 &deg;)";
      :ioos_category = "Location";
      :observation_type = "calculated";
      :platform = "platform_meta";
      :standard_name = "latitude";
      :units = "degrees_north";
      :valid_max = 90.0; // double
      :valid_min = -90.0; // double
      :references = "Rudnick, D. L., Sherman, J. T., & Wu, A. P. (2018). Depth-average velocity from Spray underwater gliders. Journal of Atmospheric and Oceanic Technology, (2018), 35, 1665-1673; doi: https://doi.org/10.1175/JTECH-D-17-0200.1";
      :accuracy = 0.007; // double
      :_ChunkSizes = 372U; // uint

    int latitude_qc(n_measurements=372);
      :_FillValue = -127; // int
      :coverage_content_type = "qualityInformation";
      :long_name = "Quality Flag for the Estimated Subsurface Latitude";
      :short_name = "Quality Flag for Subsurface Latitude";
      :standard_name = "aggregate_quality_flag";
      :valid_max = 9; // int
      :valid_min = 0; // int
      :flag_values = 1, 2, 3, 4, 9; // int
      :flag_meanings = "good not_evaluated questionable bad missing";
      :comment = "Use caution - these are estimated subsurface position values, the deviation from actual position may be several hundreds of meters! These are estimations and are a dead reckoning using the GPS positions at dive start and end, and the gliders estimated velocity. The calculation methods are described in Rudnick, D. L., Sherman, J. T., & Wu, A. P. (2018). Depth-average velocity from Spray underwater gliders. Journal of Atmospheric and Oceanic Technology, (2018), 35, 1665-1673; doi: https://doi.org/10.1175/JTECH-D-17-0200.1. The accuracy attribute reflects an accuracy of approximately +/-800m (0.09 &deg; Lon) 1=Good/Pass, 2=Not Evaluated, 3=Questionable, Suspect or of High Interest, 4=Fail/Bad, 9=Missing Data. See the references for more details on the flag meanings.";
      :references = "Paris. Intergovernmental Oceanographic Commission of UNESCO, 2013. Ocean Data Standards, Vol.3:Recommendation for a Quality Flag Scheme for the Exchange of Oceanographic and Marine    Meteorological Data. (IOC Manuals and Guides, 54, Vol. 3.) 12 pp. (English.)(IOC/2013/MG/54-3) https://repository.oceanbestpractices.org/bitstream/handle/11329/413/MG54_3.doc";
      :_ChunkSizes = 372U; // uint

    double longitude(n_measurements=372);
      :_FillValue = -999.0; // double
      :axis = "X";
      :colorBarMaximum = 180.0; // double
      :colorBarMinimum = -180.0; // double
      :comment = "Use caution - these are estimated positions of the glider underwater during a dive. Use the GPS position variables for accurate positions at the surface. Use caution with these estimated subsurface position values, the deviation from actual position may be several hundreds of meters! These estimations are a dead reckoning using the GPS positions at dive start and end, and the gliders estimated velocity. The calculation methods are described in: \'Rudnick, D. L., Sherman, J. T., & Wu, A. P. (2018). Depth-average velocity from Spray underwater gliders. Journal of Atmospheric and Oceanic Technology, (2018), 35, 1665-1673; doi: https://doi.org/10.1175/JTECH-D-17-0200.1\'. The accuracy attribute reflects an accuracy of approximately +/-800m (0.09 &deg; Lon)";
      :ioos_category = "Location";
      :long_name = "Estimated Subsurface Longitude";
      :observation_type = "calculated";
      :platform = "platform_meta";
      :standard_name = "longitude";
      :units = "degrees_east";
      :valid_max = 180.0; // double
      :valid_min = -180.0; // double
      :accuracy = 0.09; // double
      :_ChunkSizes = 372U; // uint

    int longitude_qc(n_measurements=372);
      :_FillValue = -127; // int
      :coverage_content_type = "qualityInformation";
      :long_name = "Estimated Subsurface Longitude Quality Flag";
      :standard_name = "aggregate_quality_flag";
      :valid_max = 9; // int
      :valid_min = 0; // int
      :flag_values = 1, 2, 3, 4, 9; // int
      :flag_meanings = "good not_evaluated questionable bad missing";
      :comment = "Use caution - these are estimated subsurface position values, the deviation from actual position may be several hundreds of meters! Use the gps position variables for highly accurate positions at the surface. These estimations are a dead reckoning using the GPS positions at dive start and end, and the gliders estimated velocity. The calculation methods are described in: \"Rudnick, D. L., Sherman, J. T., & Wu, A. P. (2018). Depth-average velocity from Spray underwater gliders. Journal of Atmospheric and Oceanic Technology, (2018), 35, 1665-1673; doi: https://doi.org/10.1175/JTECH-D-17-0200.1\". The accuracy attribute reflects an accuracy of approximately +/-800m (0.09 &deg; Lon)1=Good/Pass, 2=Not Evaluated, 3=Questionable, Suspect or of High Interest, 4=Fail/Bad, 9=Missing Data. See the references for more details on the flag meanings.";
      :references = "Paris. Intergovernmental Oceanographic Commission of UNESCO, 2013. Ocean Data Standards, Vol.3:Recommendation for a Quality Flag Scheme for the Exchange of Oceanographic and Marine    Meteorological Data. (IOC Manuals and Guides, 54, Vol. 3.) 12 pp. (English.)(IOC/2013/MG/54-3) https://repository.oceanbestpractices.org/bitstream/handle/11329/413/MG54_3.doc";
      :_ChunkSizes = 372U; // uint

    double pres(n_measurements=372);
      :_FillValue = -999.0; // double
      :ancillary_variables = "pres_qc";
      :coordinates = "time longitude latitude depth";
      :coverage_content_type = "physicalMeasurement";
      :long_name = "Pressure";
      :observation_type = "measured";
      :platform = "platform_meta";
      :positive = "down";
      :reference_datum = "sea-surface";
      :sensor = "sensor_ctd";
      :standard_name = "sea_water_pressure";
      :units = "dbar";
      :valid_max = 2000.0; // double
      :valid_min = 0.0; // double
      :vocabulary = "https://vocab.nerc.ac.uk/collection/OG1/current";
      :_ChunkSizes = 372U; // uint

    int pres_qc(n_measurements=372);
      :_FillValue = -127; // int
      :coordinates = "time longitude latitude depth";
      :coverage_content_type = "qualityInformation";
      :long_name = "Pressure Quality Flag";
      :standard_name = "aggregate_quality_flag";
      :valid_max = 9; // int
      :valid_min = 0; // int
      :flag_values = 1, 2, 3, 4, 9; // int
      :flag_meanings = "good not_evaluated questionable bad missing";
      :comment = "1=Good/Pass, 2=Not Evaluated, 3=Questionable, Suspect or of High Interest, 4=Fail/Bad, 9=Missing Data. See the references for more details on the flag meanings.";
      :references = "Paris. Intergovernmental Oceanographic Commission of UNESCO, 2013. Ocean Data Standards, Vol.3:Recommendation for a Quality Flag Scheme for the Exchange of Oceanographic and Marine    Meteorological Data. (IOC Manuals and Guides, 54, Vol. 3.) 12 pp. (English.)(IOC/2013/MG/54-3) https://repository.oceanbestpractices.org/bitstream/handle/11329/413/MG54_3.doc";
      :_ChunkSizes = 372U; // uint

    double psal(n_measurements=372);
      :_FillValue = -999.0; // double
      :ancillary_variables = "psal_qc";
      :colorBarMaximum = 35.0; // double
      :colorBarMinimum = 32.0; // double
      :comment = "PSS-78, calculated on board glider";
      :coordinates = "time longitude latitude depth";
      :coverage_content_type = "physicalMeasurement";
      :ioos_category = "Salinity";
      :long_name = "Sea Water Practical Salinity";
      :observation_type = "measured";
      :sensor = "sensor_ctd";
      :standard_name = "sea_water_practical_salinity";
      :units = "1";
      :valid_max = 40.0; // double
      :valid_min = 0.0; // double
      :vocabulary = "https://vocab.nerc.ac.uk/collection/OG1/current";
      :_ChunkSizes = 372U; // uint

    int psal_qc(n_measurements=372);
      :_FillValue = -127; // int
      :coverage_content_type = "qualityInformation";
      :long_name = "Sea Water Practical Salinity Quality Flag";
      :short_name = "Salinity Quality Flag";
      :valid_max = 9; // int
      :valid_min = 1; // int
      :flag_values = 1, 2, 3, 4, 9; // int
      :flag_meanings = "good not_evaluated questionable bad missing";
      :comment = "1=Good/Pass, 2=Not Evaluated, 3=Questionable, Suspect or of High Interest, 4=Fail/Bad, 9=Missing Data. See the references for more details on the flag meanings.";
      :references = "Paris. Intergovernmental Oceanographic Commission of UNESCO, 2013. Ocean Data Standards, Vol.3:Recommendation for a Quality Flag Scheme for the Exchange of Oceanographic and Marine    Meteorological Data. (IOC Manuals and Guides, 54, Vol. 3.) 12 pp. (English.)(IOC/2013/MG/54-3) https://repository.oceanbestpractices.org/bitstream/handle/11329/413/MG54_3.doc";
      :_ChunkSizes = 372U; // uint

    double temp(n_measurements=372);
      :_FillValue = -999.0; // double
      :ancillary_variables = "temp_qc";
      :colorBarMaximum = 32.0; // double
      :colorBarMinimum = 0.0; // double
      :coordinates = "time longitude latitude depth";
      :coverage_content_type = "physicalMeasurement";
      :ioos_category = "Temperature";
      :long_name = "Sea Water Temperature";
      :sensor = "sensor_ctd";
      :observation_type = "measured";
      :standard_name = "sea_water_temperature";
      :units = "degree_C";
      :valid_max = 40.0; // double
      :valid_min = -5.0; // double
      :vocabulary = "https://vocab.nerc.ac.uk/collection/OG1/current";
      :_ChunkSizes = 372U; // uint

    int temp_qc(n_measurements=372);
      :_FillValue = -127; // int
      :coordinates = "time longitude latitude depth";
      :coverage_content_type = "qualityInformation";
      :long_name = "Sea Water Temperature Quality Flag";
      :valid_max = 9; // int
      :valid_min = 1; // int
      :flag_values = 1, 2, 3, 4, 9; // int
      :flag_meanings = "good not_evaluated questionable bad missing";
      :comment = "1=Good/Pass, 2=Not Evaluated, 3=Questionable, Suspect or of High Interest, 4=Fail/Bad, 9=Missing Data. See the references for more details on the flag meanings.";
      :references = "Paris. Intergovernmental Oceanographic Commission of UNESCO, 2013. Ocean Data Standards, Vol.3:Recommendation for a Quality Flag Scheme for the Exchange of Oceanographic and Marine    Meteorological Data. (IOC Manuals and Guides, 54, Vol. 3.) 12 pp. (English.)(IOC/2013/MG/54-3) https://repository.oceanbestpractices.org/bitstream/handle/11329/413/MG54_3.doc";
      :_ChunkSizes = 372U; // uint

    double cndc(n_measurements=372);
      :_FillValue = -999.0; // double
      :ancillary_variables = "psal_qc";
      :colorBarMaximum = 6.0; // double
      :colorBarMinimum = 2.0; // double
      :coordinates = "time longitude latitude depth";
      :coverage_content_type = "physicalMeasurement";
      :long_name = "Conductivity";
      :sensor = "sensor_ctd";
      :standard_name = "sea_water_electrical_conductivity";
      :ioos_category = "salinity";
      :observation_type = "calculated";
      :platform = "platform_meta";
      :units = "S m-1";
      :valid_max = 10.0; // double
      :valid_min = 0.0; // double
      :vocabulary = "https://vocab.nerc.ac.uk/collection/OG1/current";
      :_ChunkSizes = 372U; // uint

    int cndc_qc(n_measurements=372);
      :_FillValue = -127; // int
      :comment = "1=Good/Pass, 2=Not Evaluated, 3=Questionable, Suspect or of High Interest, 4=Fail/Bad, 9=Missing Data. See the references for more details on the flag meanings.";
      :coverage_content_type = "qualityInformation";
      :long_name = "Conductivity Quality Flag";
      :valid_max = 9; // int
      :valid_min = 1; // int
      :flag_values = 1, 2, 3, 4, 9; // int
      :flag_meanings = "good not_evaluated questionable bad missing";
      :references = "Paris. Intergovernmental Oceanographic Commission of UNESCO, 2013. Ocean Data Standards, Vol.3:Recommendation for a Quality Flag Scheme for the Exchange of Oceanographic and Marine    Meteorological Data. (IOC Manuals and Guides, 54, Vol. 3.) 12 pp. (English.)(IOC/2013/MG/54-3) https://repository.oceanbestpractices.org/bitstream/handle/11329/413/MG54_3.doc";
      :_ChunkSizes = 372U; // uint

    double chla(n_measurements=372);
      :_FillValue = -999.0; // double
      :ancillary_variables = "chla_qc";
      :comment = "Chlorophyll-a concentration estimated from fluorescence measurements. See the sensor_fchl variable for information about the fluorometer.";
      :coordinates = "time longitude latitude depth";
      :coverage_content_type = "physicalMeasurement";
      :ioos_category = "Other";
      :long_name = "Chlorophyll-a concentration";
      :observation_type = "measured";
      :sensor = "sensor_fchl";
      :standard_name = "mass_concentration_of_chlorophyll_a_in_sea_water";
      :units = "mg m-3";
      :vocabulary = "https://vocab.nerc.ac.uk/collection/OG1/current";
      :_ChunkSizes = 372U; // uint

    int chla_qc(n_measurements=372);
      :_FillValue = -127; // int
      :coordinates = "time longitude latitude depth";
      :coverage_content_type = "qualityInformation";
      :long_name = "Chlorophyll-a concentration Quality Flag";
      :valid_max = 9; // int
      :valid_min = 1; // int
      :flag_values = 1, 2, 3, 4, 9; // int
      :flag_meanings = "good not_evaluated questionable bad missing";
      :comment = "1=Good/Pass, 2=Not Evaluated, 3=Questionable, Suspect or of High Interest, 4=Fail/Bad, 9=Missing Data. See the references for more details on the flag meanings.";
      :references = "Paris. Intergovernmental Oceanographic Commission of UNESCO, 2013. Ocean Data Standards, Vol.3:Recommendation for a Quality Flag Scheme for the Exchange of Oceanographic and Marine    Meteorological Data. (IOC Manuals and Guides, 54, Vol. 3.) 12 pp. (English.)(IOC/2013/MG/54-3) https://repository.oceanbestpractices.org/bitstream/handle/11329/413/MG54_3.doc";
      :_ChunkSizes = 372U; // uint

    double doxy(n_measurements=372);
      :_FillValue = -999.0; // double
      :ancillary_variables = "doxy_qc";
      :coordinates = "time longitude latitude depth";
      :coverage_content_type = "physicalMeasurement";
      :ioos_category = "physical_oceanography";
      :long_name = "Dissolved Oxygen";
      :observation_type = "measured";
      :platform = "platform_meta";
      :sensor = "sensor_doxy";
      :standard_name = "moles_of_oxygen_per_unit_mass_in_sea_water";
      :units = "micromol kg-1";
      :valid_max = 500.0; // double
      :valid_min = 0.0; // double
      :vocabulary = "https://vocab.nerc.ac.uk/collection/OG1/current";
      :_ChunkSizes = 372U; // uint

    int doxy_qc(n_measurements=372);
      :_FillValue = -127; // int
      :coordinates = "time longitude latitude depth";
      :coverage_content_type = "qualityInformation";
      :long_name = "Dissolved Oxygen Quality Flag";
      :valid_max = 9; // int
      :valid_min = 1; // int
      :flag_values = 1, 2, 3, 4, 9; // int
      :flag_meanings = "good not_evaluated questionable bad missing";
      :comment = "1=Good/Pass, 2=Not Evaluated, 3=Questionable, Suspect or of High Interest, 4=Fail/Bad, 9=Missing Data. See the references for more details on the flag meanings.";
      :references = "Paris. Intergovernmental Oceanographic Commission of UNESCO, 2013. Ocean Data Standards, Vol.3:Recommendation for a Quality Flag Scheme for the Exchange of Oceanographic and Marine    Meteorological Data. (IOC Manuals and Guides, 54, Vol. 3.) 12 pp. (English.)(IOC/2013/MG/54-3) https://repository.oceanbestpractices.org/bitstream/handle/11329/413/MG54_3.doc";
      :_ChunkSizes = 372U; // uint

    double time_gps(n_measurements=372);
      :_FillValue = -999.0; // double
      :ancillary_variables = "gps_start_qc gps_start_qc_tests";
      :calendar = "gregorian";
      :comment = "Time from GPS at surface for the start position of the dive. These data are transmitted in near-real-time and are uncorrected. Flags are provided in the gps_start_qc and gps_start_qc_tests variables. ";
      :ioos_category = "Time";
      :long_name = "GPS Time at Dive Start";
      :observation_type = "measured";
      :platform = "platform_meta";
      :standard_name = "time";
      :units = "seconds since 1970-01-01T00:00:00Z";
      :valid_min = 1.0E9; // double
      :valid_max = 4.0E9; // double
      :_ChunkSizes = 372U; // uint

    double longitude_gps(n_measurements=372);
      :_FillValue = -999.0; // double
      :_CoordinateAxisType = "Lon";
      :ancillary_variables = "gps_start_qc gps_start_qc_tests";
      :comment = "Longitude from GPS at surface for the starting position of the dive. These data are transmitted in near-real-time and are uncorrected. Flags are provided in the gps_end_qc and gps_end_qc_tests variables. ";
      :ioos_category = "Location";
      :long_name = "GPS Longitude at Dive Start";
      :observation_type = "measured";
      :platform = "platform_meta";
      :standard_name = "longitude";
      :units = "degrees_east";
      :valid_max = 180.0; // double
      :valid_min = -180.0; // double
      :_ChunkSizes = 372U; // uint

    double latitude_gps(n_measurements=372);
      :_FillValue = -999.0; // double
      :ancillary_variables = "gps_start_qc gps_start_qc_tests";
      :comment = "Latitude from GPS at surface for the start position of the dive. These data are transmitted in near-real-time and are uncorrected. Flags are provided in the gps_start_qc and gps_start_qc_tests variables. ";
      :ioos_category = "Location";
      :long_name = "GPS Latitude at Dive Start";
      :observation_type = "measured";
      :platform = "platform_meta";
      :standard_name = "latitude";
      :units = "degrees_north";
      :valid_max = 90.0; // double
      :valid_min = -90.0; // double
      :_ChunkSizes = 372U; // uint

    int gps_start_qc(n_measurements=372);
      :_FillValue = -127; // int
      :comment = "1=Good/Pass, 2=Not Evaluated, 3=Questionable, Suspect or of High Interest, 4=Fail/Bad, 9=Missing Data. See the references for more details on the flag meanings.";
      :flag_values = 1, 2, 3, 4, 9; // int
      :flag_meanings = "good not_evaluated questionable bad missing";
      :long_name = "Summary Quality Flag for the GPS Start Position";
      :references = "Paris. Intergovernmental Oceanographic Commission of UNESCO, 2013. Ocean Data Standards, Vol.3:Recommendation for a Quality Flag Scheme for the Exchange of Oceanographic and Marine    Meteorological Data. (IOC Manuals and Guides, 54, Vol. 3.) 12 pp. (English.)(IOC/2013/MG/54-3) https://repository.oceanbestpractices.org/bitstream/handle/11329/413/MG54_3.doc";
      :standard_name = "aggregate_quality_flag";
      :valid_max = 9; // int
      :valid_min = 1; // int
      :_ChunkSizes = 372U; // uint

    int gps_start_qc_tests(n_measurements=372);
      :_FillValue = -127; // int
      :comment = "gps_good=0 gps_day_problem=1 gps_repeat=2 gps_backward=3 gps_too_fast_on_surface=4 gps_too_soon=5 gps_too_far=6 gps_bad_hdop=7 gps_bad_status=8 gps_no_surfacing=9 gps_manual=10 gps_no_dive=99";
      :long_name = "Detailed Quality Flags for the GPS Start Position";
      :flag_values = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 99; // int
      :flag_meanings = "gps_good gps_day_problem gps_repeat gps_backward gps_too_fast_on_surface gps_too_soon gps_too_far gps_bad_hdop gps_bad_status gps_no_surfacing gps_manual gps_no_dive";
      :standard_name = "quality_flag";
      :valid_max = 99; // int
      :valid_min = 0; // int
      :_ChunkSizes = 372U; // uint

    double time_gps_end(n_measurements=372);
      :_FillValue = -999.0; // double
      :ancillary_variables = "gps_end_qc gps_end_qc_tests";
      :comment = "Time from GPS at surface for the end position of the dive. These data are transmitted in near-real-time. Flags are provided in the gps_start_qc and gps_start_qc_tests variables. This location corresponds closely with the surface value of the profile measurements.";
      :ioos_category = "Location";
      :long_name = "GPS Time at Dive End";
      :observation_type = "measured";
      :platform = "platform_meta";
      :standard_name = "time";
      :units = "seconds since 1970-01-01T00:00:00Z";
      :valid_min = 1.0E9; // double
      :valid_max = 4.0E9; // double
      :_ChunkSizes = 372U; // uint

    double latitude_gps_end(n_measurements=372);
      :_FillValue = -999.0; // double
      :colorBarMaximum = 90.0; // double
      :colorBarMinimum = -90.0; // double
      :comment = "Latitude from GPS at surface for the end position of the dive. These data are transmitted in near-real-time. Flags are provided in the gps_start_qc and gps_start_qc_tests variables.This location corresponds closely with the surface value of the profile measurements.";
      :ioos_category = "Location";
      :long_name = "GPS Latitude at Dive End";
      :observation_type = "measured";
      :platform = "platform_meta";
      :standard_name = "latitude";
      :units = "degrees_north";
      :valid_max = 90.0; // double
      :valid_min = -90.0; // double
      :ancillary_variables = "gps_end_qc gps_end_qc_tests";
      :_ChunkSizes = 372U; // uint

    double longitude_gps_end(n_measurements=372);
      :_FillValue = -999.0; // double
      :colorBarMaximum = 180.0; // double
      :colorBarMinimum = -180.0; // double
      :comment = "Longitude from GPS at surface for the ending position of the dive. These data are transmitted in near-real-time. Flags are provided in the gps_end_qc and gps_end_qc_tests variables. This location corresponds closely with the surface position of the profile measurements.";
      :ioos_category = "Location";
      :long_name = "GPS Longitude at Dive End";
      :observation_type = "measured";
      :platform = "platform_meta";
      :standard_name = "longitude";
      :units = "degrees_east";
      :valid_max = 180.0; // double
      :valid_min = -180.0; // double
      :ancillary_variables = "gps_end_qc gps_end_qc_tests";
      :_ChunkSizes = 372U; // uint

    int gps_end_qc(n_measurements=372);
      :_FillValue = -127; // int
      :long_name = "Summary Quality Flag for the GPS End Postion";
      :valid_max = 9; // int
      :valid_min = 1; // int
      :flag_values = 1, 2, 3, 4, 9; // int
      :flag_meanings = "good not_evaluated questionable bad missing";
      :comment = "1=Good/Pass, 2=Not Evaluated, 3=Questionable, Suspect or of High Interest, 4=Fail/Bad, 9=Missing Data. See the references for more details on the flag meanings.";
      :references = "Paris. Intergovernmental Oceanographic Commission of UNESCO, 2013. Ocean Data Standards, Vol.3:Recommendation for a Quality Flag Scheme for the Exchange of Oceanographic and Marine    Meteorological Data. (IOC Manuals and Guides, 54, Vol. 3.) 12 pp. (English.)(IOC/2013/MG/54-3) https://repository.oceanbestpractices.org/bitstream/handle/11329/413/MG54_3.doc";
      :standard_name = "aggregate_quality_flag";
      :_ChunkSizes = 372U; // uint

    int gps_end_qc_tests(n_measurements=372);
      :_FillValue = -127; // int
      :long_name = "Detailed Quality Flags for the GPS End Position";
      :valid_max = 99; // int
      :valid_min = 0; // int
      :flag_values = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 99; // int
      :flag_meanings = "gps_good gps_day_problem gps_repeat gps_backward gps_too_fast_on_surface gps_too_soon gps_too_far gps_bad_hdop gps_bad_status gps_no_surfacing gps_manual gps_no_dive";
      :comment = "gps_good=0 gps_day_problem=1 gps_repeat=2 gps_backward=3 gps_too_fast_on_surface=4 gps_too_soon=5 gps_too_far=6 gps_bad_hdop=7 gps_bad_status=8 gps_no_surfacing=9 gps_manual=10 gps_no_dive=99";
      :standard_name = "quality_flag";
      :_ChunkSizes = 372U; // uint

    String wmo_identifier;
      :ioos_category = "Identifier";
      :long_name = "WMO ID";

    int sensor_doxy;
      :_FillValue = -127; // int
      :_Unsigned = "false";
      :coverage_content_type = "referenceInformation";
      :ioos_category = "Identifier";
      :long_name = "Oxygen Sensor Metadata";
      :make_model = "Sea-Bird SBE 63 dissolved oxygen sensor";
      :platform = "platform_meta";
      :type = "OPTODE_DOXY";
      :type_vocabulary = "http://vocab.nerc.ac.uk/collection/R25/current/";
      :maker = "Sea-Bird Scientific";
      :maker_vocabulary = "http://vocab.nerc.ac.uk/collection/R26/current/";
      :model = "Sea-Bird SBE 63 dissolved oxygen sensor";
      :model_vocabulary = "http://vocab.nerc.ac.uk/collection/L22/current/";

    int sensor_ctd;
      :_FillValue = -127; // int
      :_Unsigned = "false";
      :coverage_content_type = "referenceInformation";
      :ioos_category = "Identifier";
      :long_name = "CTD Metadata";
      :make_model = "Sea-Bird SBE 41CP CTD";
      :platform = "platform_meta";
      :type = "CTD";
      :units = "1";
      :maker = "Sea-Bird Scientific";
      :maker_vocabulary = "https://vocab.nerc.ac.uk/collection/L35/current";
      :maker_uri = "https://vocab.nerc.ac.uk/collection/L35/current/MAN0013/";
      :model = "Sea-Bird SBE 41CP CTD";
      :model_vocabulary = "https://vocab.nerc.ac.uk/collection/L22/current";
      :model_uri = "https://vocab.nerc.ac.uk/collection/L22/current/TOOL0669/";
      :type_vocabulary = "https://vocab.nerc.ac.uk/collection/L05/current";
      :type_uri = "https://vocab.nerc.ac.uk/collection/L05/current/130/";

    int sensor_fchl;
      :_FillValue = -127; // int
      :_Unsigned = "false";
      :coverage_content_type = "referenceInformation";
      :ioos_category = "Identifier";
      :long_name = "Fluorometer Metadata";
      :platform = "platform_meta";
      :type = "fluorometer_chla";
      :type_vocabulary = "http://vocab.nerc.ac.uk/collection/R25/current/";
      :maker = "Seapoint Sensors, Inc.";
      :maker_vocabulary = "http://vocab.nerc.ac.uk/collection/R26/current/";
      :model = "Seapoint chlorophyll fluorometer";
      :model_vocabulary = "http://vocab.nerc.ac.uk/collection/L05/current";
      :model_uri = "http://vocab.nerc.ac.uk/collection/L05/current/113/";

    String platform_model;
      :ioos_category = "Identifier";
      :long_name = "Model of the glider";
      :comment = "The NERC vocabulary defines terms used to describe designs or versions of platforms.";
      :platform_model_uri = "http://vocab.nerc.ac.uk/collection/B76/current/B7600027/";
      :platform_model_vocabulary = "http://vocab.nerc.ac.uk/collection/B76/current/";

    String platform_serial_number;
      :ioos_category = "Identifier";
      :long_name = "Glider serial number";

    int platform_meta;
      :_FillValue = -127; // int
      :comment = "Spray Glider sp028";
      :coverage_content_type = "referenceInformation";
      :id = "sp028";
      :sensor = "sensor_ctd";
      :ioos_category = "Identifier";
      :long_name = "Platform Metadata";
      :platform_type = "subsurface gliders";
      :platform_type_vocabulary = "http://vocab.nerc.ac.uk/collection/L06/current/27/";
      :platform_maker = "Scripps Institution of Oceanography Instrument Development Group";
      :platform_depth_rating = "1000";
      :platform_model = "Scripps Institution of Oceanography Spray glider";
      :platform_model_uri = "http://vocab.nerc.ac.uk/collection/B76/current/B7600027/";
      :platform_model_vocabulary = "http://vocab.nerc.ac.uk/collection/B76/current/";
      :platform_serial_number = "sp028";
      :type = "platform";
      :units = "1";
      :wmo_id = "4801921";
      :wmo_identifier = "4801921";

    double deployment_time(n_measurements=372);
      :_FillValue = -999.0; // double
      :comment = "GPS Time value for the start position of the first dive.";
      :ioos_category = "Location";
      :long_name = "Deployment Time, GPS at start of first dive";
      :observation_type = "measured";
      :platform = "platform_meta";
      :standard_name = "time";
      :units = "seconds since 1970-01-01T00:00:00Z";
      :_ChunkSizes = 372U; // uint

    double deployment_latitude(n_measurements=372);
      :_FillValue = -999.0; // double
      :comment = "GPS latitude value for the start position of the first dive.";
      :ioos_category = "Location";
      :long_name = "Deployment Latitude, GPS at start of first dive";
      :observation_type = "measured";
      :platform = "platform_meta";
      :standard_name = "latitude";
      :units = "degrees_north";
      :_ChunkSizes = 372U; // uint

    double deployment_longitude(n_measurements=372);
      :_FillValue = -999.0; // double
      :comment = "GPS longitude value for the start position of the first dive.";
      :ioos_category = "Location";
      :long_name = "Deployment longitude, GPS at start of first dive";
      :observation_type = "measured";
      :platform = "platform_meta";
      :standard_name = "longitude";
      :units = "degrees_east";
      :_ChunkSizes = 372U; // uint

  // global attributes:
  :Conventions = "CF-1.10, ACDD-1.3, OG-1.0";
  :acknowledgement = "Funded by National Oceanic and Atmospheric Administration (NOAA): Global Ocean Monitoring and Observing (GOMO) Program and Integrated Ocean Observing System. Supported by Instrument Development Group - Scripps Institution of Oceanography";
  :cdm_trajectory_variables = "trajectory";
  :comment = "CAUTION! This is an experimental truncated file to be used solely as an OG-1.0 format example. Visit the U.S. Glider DAC at https://gliders.ioos.us/erddap/info/sp028-20230202T1637/index.html to view the NRT data. This file contains data from the following specific sensors: Sea-Bird SBE 41CP CTD, Seapoint chlorophyll fluorometer, Sea-Bird SBE 63 dissolved oxygen sensor.";
  :contributing_institutions = "Scripps Institution of Oceanography";
  :contributing_institutions_role = "Operator";
  :contributing_institutions_vocabulary = "https://vocab.nerc.ac.uk/collection/W08/current/";
  :contributor_email = "drudnick@ucsd.edu, jpsevadjian@ucsd.edu";
  :contributor_name = "Daniel Rudnick, Jennifer Sevadjian";
  :contributor_role = "principalInvestigator, resourceProvider";
  :contributor_role_vocabulary = "https://vocab.nerc.ac.uk/collection/G04/current";
  :creator_email = "idgdata@ucsd.edu";
  :creator_institution = "Scripps Institution of Oceanography";
  :creator_name = "Instrument Development Group";
  :creator_type = "group";
  :creator_url = "https://spraydata.ucsd.edu";
  :data_url = "https://spraydata.ucsd.edu/erddap/info/sp028_20230202T1637_R/index.html";
  :date_created = "2024-06-07T19:40:02Z";
  :date_issued = "2024-06-07T19:40:02Z";
  :date_metadata_modified = "2024-06-07T19:40:02Z";
  :date_modified = "2024-06-07T19:40:02Z";
  :doi = "10.21238/S8SPRAY1618";
  :featureType = "trajectory";
  :geospatial_bounds = "POLYGON ((-123.36765 38.318775, -123.0713 38.318775, -123.0713 38.246275, -123.36765 38.246275, -123.36765 38.318775))";
  :geospatial_bounds_crs = "EPSG:4326";
  :geospatial_lat_max = 38.318775; // double
  :geospatial_lat_min = 38.246275; // double
  :geospatial_lat_units = "degrees_north";
  :geospatial_lon_max = -123.0713; // double
  :geospatial_lon_min = -123.36765; // double
  :geospatial_lon_units = "degrees_east";
  :geospatial_vertical_max = 0.03969955209296338; // double
  :geospatial_vertical_min = 111.36731572605271; // double
  :geospatial_vertical_positive = "down";
  :geospatial_vertical_units = "EPSG:5831";
  :history = "2023-06-16T15:40:09Z: Jenn readsat(maxdives=3000, Gps_Good=0, Gps_Bad=8, Gps_No_Dive=99, Gps_No_Surfacing=9, DOConv=44660). \n2023-06-16T15:40:49Z: Jenn fixgps3(R=6378000, Too_Soon=60, Too_Fast_On_Surface=5, Too_Far=100, Bad_HDOP=12, Gps_Good=0, Gps_Repeat=2, Gps_Backward=3, Gps_Too_Fast_On_Surface=4, Gps_Too_Soon=5, Gps_Too_Far=6, Gps_Bad_HDOP=7, Gps_Bad_Status=8, Gps_No_Surfacing=9). \n2023-06-16T15:40:49Z: Jenn calcvelsat(R=6378000, Gps_No_Surfacing=9). \n2023-06-16T15:42:15Z: Jenn calox(filename=/Users/Shared/spray/data/ox/doxcal.xlsx, sheetname=AllOxMissions, DOConv=44660, Gain=1.0811, Offset=-0.0615). \n;2024-06-07T19:40:02Z: OG-1.0 NetCDF created by J.P. Sevadjian with make_mission_nc_og10.py, input file: 23202801_aug.mat, with MD5 checksum: b0936e175fd11895c04fdba38f379df0, output file: ./mission_output/OG-10-202400415/20240607/sp028_20230202T1637_R.nc.";
  :id = "sp028_20230202T1637";
  :infoUrl = "https://spraydata.ucsd.edu";
  :institution = "Scripps Institution of Oceanography";
  :instrument = "CAUTION! This is an experimental truncated file to be used solely as an OG-1.0 format example. Visit the U.S. Glider DAC at https://gliders.ioos.us/erddap/info/sp028-20230202T1637/index.html to view the NRT data. This file contains data from the following specific sensors: Sea-Bird SBE 41CP CTD, Seapoint chlorophyll fluorometer, Sea-Bird SBE 63 dissolved oxygen sensor.";
  :internal_mission_identifier = "23202801";
  :keywords = "AUVS > Autonomous Underwater Vehicles, Earth Science > Oceans > Ocean Pressure > Water Pressure, Earth Science > Oceans > Ocean Temperature > Water Temperature, Earth Science > Oceans > Salinity/Density > Conductivity, Earth Science > Oceans > Salinity/Density > Density, Earth Science > Oceans > Salinity/Density > Salinity, glider, In Situ Ocean-based platforms > Seaglider, Slocum, Spray, trajectory, underwater glider, water, wmo, underwater glider, pressure, temperature, salinity, currents, oxygen, fluorescence, chlorophyll;";
  :keywords_vocabulary = "GCMD Science Keywords";
  :license = "The data may be used and redistributed for free but is not intended for legal use, since it may contain inaccuracies. Neither the data Contributor, University of California, IOOS, NOAA, nor the United States Government, nor any of their employees or contractors, makes any warranty, express or implied, including warranties of merchantability and fitness for a particular purpose, or assumes any legal liability for the accuracy, completeness, or usefulness, of this information.";
  :metadata_link = "https://spraydata.ucsd.edu";
  :naming_authority = "edu.ucsd.idg";
  :network = "OceanGliders > BOON > Northeast Pacific Ocean > California Underwater Glider Network, California Underwater Glider Network (CUGN), IOOS";
  :platform = "sub-surface gliders";
  :platform_institution = "Scripps Institution of Oceanography";
  :platform_type = "Spray Glider";
  :platform_vocabulary = "https://vocab.nerc.ac.uk/collection/L06/current/";
  :processing_level = "This is a near-real-time data product. Within the Spray program to is considered a Level 2 product. Real-time quality control has been conducted and users should apply the supplied QARTOD flags. Afer a mission is complete a higher-quality data product is provided at https://spraydata.ucsd.edu and should be used in place of the near-real-time data as soon as it is available.";
  :project = "California Underwater Glider Network (CUGN)";
  :publisher_email = "idgdata@ucsd.edu";
  :publisher_institution = "University of California - San Diego; Scripps Institution of Oceanography";
  :publisher_name = "Instrument Development Group";
  :publisher_type = "group";
  :publisher_url = "https://spraydata.ucsd.edu";
  :references = "Rudnick, D. L. (2016). Ocean research enabled by underwater gliders. Annual review of marine science, 8, 519-541, doi:10.1146/annurev-marine-122414-033913\n Rudnick, D. L., Davis, R. E., & Sherman, J. T. (2016). Spray Underwater Glider Operations. Journal of Atmospheric and Oceanic Technology, 33(6), 1113-1122, doi:10.1175/JTECH-D-15-0252.1\n Rudnick, D. L., Davis, R. E., Eriksen, C. C., Fratantoni, D. M., & Perry, M. J. (2004). Underwater gliders for ocean research. Marine Technology Society Journal, 38(2), 73-84, doi:10.4031/002533204787522703\n Sherman, J., Davis, R. E., Owens, W. B., & Valdes, J. (2001). The autonomous underwater glider \'Spray\'. IEEE Journal of oceanic Engineering, 26(4), 437-446, doi:10.1109/48.972076";
  :rtqc_method = "Spray Data Center RTQC";
  :sea_name = "Coastal Waters of California";
  :site = "CUGN Line 56";
  :source = "Spray Underwater Glider";
  :standard_name_vocabulary = "CF Standard Name Table v83";
  :summary = "CAUTION! This is an experimental truncated file to be used solely as an OG-1.0 format example. Visit the U.S. Glider DAC at https://gliders.ioos.us/erddap/info/sp028-20230202T1637/index.html to view the NRT data. Spray glider data from mission 23202801, part of the California Underwater Glider Network (CUGN) project. This is the near-real-time dataset for the full mission, spanning from 2023-02-02 to 2023-05-25. \n\nThe overarching goal of the California Underwater Glider Network is to sustain baseline observations of climate variability off the coast of California. The technical approach is to deploy autonomous underwater gliders in a network to provide real-time data.\nThe CUGN uses Spray underwater gliders making repeated dives from the surface to 500 m and back, repeating the cycle every 3 hours, and traveling 3 km in the horizontal during that time. The CUGN includes gliders on three of the traditional cross-shore CalCOFI lines: line 66.7 off Monterey Bay, line 80 off Point Conception, and line 90 off Dana Point.\n The glider missions typically last about 100 days, and cover over 2000 km, thus providing 4-6 sections on lines extending 300-500 km offshore. Since 2005 the CUGN has covered 200,000 km over ground in 28 glider-years, while doing 90,000 dives.";
  :time_coverage_duration = "P0000-03-22T21:25:00";
  :time_coverage_end = "2023-05-25T14:02:00Z";
  :time_coverage_resolution = "P0000-00-00T00:00:04";
  :time_coverage_start = "2023-02-02T16:37:00Z";
  :title = "Example OG-1.0 Format with truncated data from Spray Glider Mission 23202801 (sp028_20230202T1637)";

  data:
    trajectory =   "sp028_20230202T1637"
    profile_index = 
      {2, 3, 4, 5, 6, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35}
    time_profile = 
      {1.675361294999998E9, 1.6753642950000005E9, 1.6753672950000026E9, 1.6753702949999971E9, 1.675373415E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9}
    time_profile_qc = 
      {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
    latitude_profile = 
      {38.3187, 38.3187, 38.318775, 38.3187, 38.3187, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275}
    latitude_profile_qc = 
      {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
    latitude_uv = 
      {38.3187, 38.3187, 38.31875, 38.3187, 38.3187, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685}
    latitude_uv_qc = 
      {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
    longitude_profile = 
      {-123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765}
    longitude_profile_qc = 
      {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
    longitude_uv = 
      {-123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366}
    longitude_uv_qc = 
      {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
    time_uv = 
      {1.6753605899999974E9, 1.6753635899999995E9, 1.675366590000002E9, 1.675369589999999E9, 1.6753727099999993E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9}
    time_uv_qc = 
      {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
    time = 
      {1.675361294999998E9, 1.6753642950000005E9, 1.6753672950000026E9, 1.6753702949999971E9, 1.675373415E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9}
    time_qc = 
      {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
    wcur_x = 
      {0.0011, 7.0E-4, 0.0011, 0.0014, 0.0011, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242}
    wcur_y = 
      {7.0E-4, 4.0E-4, 0.0043, 7.0E-4, 7.0E-4, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603}
    wcur_qc = 
      {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
    wcur_qc_tests = 
      {0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0}
    depth = 
      {0.0397, 0.0794, 0.0794, 0.0397, 0.0397, 111.3673, 111.0896, 110.3754, 109.9786, 109.066, 108.4708, 107.5979, 106.8836, 105.8916, 105.3361, 104.0664, 103.2728, 102.2411, 101.4078, 100.1778, 99.3445, 97.4398, 96.0906, 94.305, 92.8764, 91.6066, 90.2177, 88.9479, 87.6384, 85.8923, 84.5828, 83.3923, 81.9637, 80.6144, 79.5032, 78.1143, 76.9634, 75.8919, 74.5426, 73.3918, 72.3599, 70.9312, 69.701, 68.7088, 67.5579, 65.9704, 64.8195, 63.7876, 62.5176, 61.4461, 60.4935, 59.3029, 58.271, 57.3582, 56.4056, 55.1356, 54.064, 53.1511, 51.9604, 50.5713, 49.4203, 48.428, 47.0785, 46.0069, 45.0146, 43.943, 42.4744, 41.2042, 40.1326, 38.267, 36.9969, 35.8458, 34.2977, 32.9482, 31.8764, 30.3284, 29.1376, 27.9864, 26.5574, 25.4063, 24.3345, 23.0246, 21.9528, 21.0001, 19.6108, 18.4596, 17.229, 16.1572, 14.8075, 13.696, 12.8226, 11.7111, 10.7187, 9.2101, 8.1383, 6.9473, 5.9946, 5.0815, 3.8111, 2.9378, 1.9056, 108.5105, 108.1137, 107.3201, 106.5662, 105.7726, 105.0584, 104.3442, 103.3522, 102.5586, 101.6856, 100.7333, 99.781, 98.9477, 97.8366, 96.924, 95.8922, 94.9399, 93.2336, 92.0431, 90.4558, 89.2257, 88.0352, 86.8447, 85.6542, 84.305, 83.1145, 81.4478, 80.0588, 78.8286, 77.1222, 75.7729, 73.9474, 72.6774, 71.3281, 69.7407, 68.3119, 67.161, 65.4942, 64.1448, 62.9939, 61.5254, 60.2951, 59.2632, 57.8741, 56.8025, 55.8103, 54.5799, 53.5083, 52.6352, 51.3254, 50.2141, 49.1821, 48.0311, 46.6816, 45.4115, 44.2605, 42.6728, 41.3233, 40.2119, 38.6639, 37.3144, 36.0442, 34.4168, 33.0276, 31.9161, 30.2093, 28.9391, 27.9071, 26.4384, 25.2475, 24.2551, 22.8658, 21.7146, 20.6825, 19.3329, 18.142, 17.0702, 15.8396, 14.3708, 13.2196, 12.1081, 10.4805, 9.3689, 7.9398, 6.5901, 5.3991, 4.4066, 3.0172, 1.8659, 110.6531, 110.3754, 109.8199, 109.2644, 108.7089, 107.9947, 107.3995, 106.6059, 105.8917, 105.1775, 104.2648, 103.3919, 102.5586, 101.5269, 100.5746, 99.5826, 98.6302, 96.6065, 95.297, 93.5511, 92.1225, 90.9717, 89.5035, 88.3924, 87.0035, 85.1781, 83.9082, 82.678, 81.17, 79.8207, 78.6699, 77.2016, 75.892, 74.7411, 73.1537, 71.725, 70.4947, 68.6295, 67.2007, 65.2561, 63.7083, 62.4383, 60.6523, 59.2632, 57.6757, 56.3263, 55.1753, 53.7465, 52.4367, 51.2857, 49.8569, 48.6265, 47.4755, 45.9275, 44.578, 43.3873, 41.7996, 40.4898, 39.4181, 37.9495, 36.8381, 35.687, 34.1787, 33.0276, 31.8765, 30.3681, 29.1773, 27.9071, 26.5971, 25.0887, 23.8979, 22.3895, 21.1589, 20.0871, 18.7771, 17.626, 16.6335, 15.4029, 14.0532, 12.8226, 11.7508, 10.0835, 8.5353, 7.3443, 6.1137, 4.9624, 3.9699, 2.6599, 1.5086, 108.4312, 108.0741, 107.4392, 106.844, 106.0504, 105.4156, 104.5823, 103.9077, 103.1538, 102.3205, 101.4476, 100.6143, 99.7413, 98.8287, 97.797, 96.924, 95.8129, 94.2257, 93.1543, 91.7257, 90.6543, 89.6622, 88.5511, 87.5591, 86.4083, 85.2971, 84.0273, 82.6383, 81.4081, 80.2176, 78.7493, 77.4397, 76.2888, 74.3442, 72.9553, 71.2488, 69.8994, 68.6692, 67.042, 65.653, 64.4623, 62.6764, 61.327, 60.057, 58.5092, 57.1201, 55.8897, 54.3021, 52.8733, 51.3651, 50.0553, 48.8646, 47.3564, 46.1657, 45.1337, 43.4667, 42.3553, 41.2836, 39.9341, 38.8227, 37.8304, 36.719, 35.4489, 34.3772, 33.4642, 32.0352, 30.8841, 29.8521, 28.8597, 27.4704, 26.359, 25.3666, 24.0964, 22.9849, 22.0322, 20.9207, 19.7299, 18.6581, 17.7054, 16.4351, 15.3236, 14.212, 13.2196, 11.9096, 10.7981, 9.885, 7.4237, 6.4313, 5.3594, 4.089, 3.0569, 2.0644, 1.0322}
    depth_qc = 
      {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
    latitude = 
      {38.3187, 38.3187, 38.318775, 38.3187, 38.3187, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275}
    latitude_qc = 
      {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
    longitude = 
      {-123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765}
    longitude_qc = 
      {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
    pres = 
      {0.04, 0.08, 0.08, 0.04, 0.04, 112.24, 111.96, 111.24, 110.84, 109.92, 109.32, 108.44, 107.72, 106.72, 106.16, 104.88, 104.08, 103.04, 102.2, 100.96, 100.12, 98.2, 96.84, 95.04, 93.6, 92.32, 90.92, 89.64, 88.32, 86.56, 85.24, 84.04, 82.6, 81.24, 80.12, 78.72, 77.56, 76.48, 75.12, 73.96, 72.92, 71.48, 70.24, 69.24, 68.08, 66.48, 65.32, 64.28, 63.0, 61.92, 60.96, 59.76, 58.72, 57.8, 56.84, 55.56, 54.48, 53.56, 52.36, 50.96, 49.8, 48.8, 47.44, 46.36, 45.36, 44.28, 42.8, 41.52, 40.44, 38.56, 37.28, 36.12, 34.56, 33.2, 32.12, 30.56, 29.36, 28.2, 26.76, 25.6, 24.52, 23.2, 22.12, 21.16, 19.76, 18.6, 17.36, 16.28, 14.92, 13.8, 12.92, 11.8, 10.8, 9.28, 8.2, 7.0, 6.04, 5.12, 3.84, 2.96, 1.92, 109.36, 108.96, 108.16, 107.4, 106.6, 105.88, 105.16, 104.16, 103.36, 102.48, 101.52, 100.56, 99.72, 98.6, 97.68, 96.64, 95.68, 93.96, 92.76, 91.16, 89.92, 88.72, 87.52, 86.32, 84.96, 83.76, 82.08, 80.68, 79.44, 77.72, 76.36, 74.52, 73.24, 71.88, 70.28, 68.84, 67.68, 66.0, 64.64, 63.48, 62.0, 60.76, 59.72, 58.32, 57.24, 56.24, 55.0, 53.92, 53.04, 51.72, 50.6, 49.56, 48.4, 47.04, 45.76, 44.6, 43.0, 41.64, 40.52, 38.96, 37.6, 36.32, 34.68, 33.28, 32.16, 30.44, 29.16, 28.12, 26.64, 25.44, 24.44, 23.04, 21.88, 20.84, 19.48, 18.28, 17.2, 15.96, 14.48, 13.32, 12.2, 10.56, 9.44, 8.0, 6.64, 5.44, 4.44, 3.04, 1.88, 111.52, 111.24, 110.68, 110.12, 109.56, 108.84, 108.24, 107.44, 106.72, 106.0, 105.08, 104.2, 103.36, 102.32, 101.36, 100.36, 99.4, 97.36, 96.04, 94.28, 92.84, 91.68, 90.2, 89.08, 87.68, 85.84, 84.56, 83.32, 81.8, 80.44, 79.28, 77.8, 76.48, 75.32, 73.72, 72.28, 71.04, 69.16, 67.72, 65.76, 64.2, 62.92, 61.12, 59.72, 58.12, 56.76, 55.6, 54.16, 52.84, 51.68, 50.24, 49.0, 47.84, 46.28, 44.92, 43.72, 42.12, 40.8, 39.72, 38.24, 37.12, 35.96, 34.44, 33.28, 32.12, 30.6, 29.4, 28.12, 26.8, 25.28, 24.08, 22.56, 21.32, 20.24, 18.92, 17.76, 16.76, 15.52, 14.16, 12.92, 11.84, 10.16, 8.6, 7.4, 6.16, 5.0, 4.0, 2.68, 1.52, 109.28, 108.92, 108.28, 107.68, 106.88, 106.24, 105.4, 104.72, 103.96, 103.12, 102.24, 101.4, 100.52, 99.6, 98.56, 97.68, 96.56, 94.96, 93.88, 92.44, 91.36, 90.36, 89.24, 88.24, 87.08, 85.96, 84.68, 83.28, 82.04, 80.84, 79.36, 78.04, 76.88, 74.92, 73.52, 71.8, 70.44, 69.2, 67.56, 66.16, 64.96, 63.16, 61.8, 60.52, 58.96, 57.56, 56.32, 54.72, 53.28, 51.76, 50.44, 49.24, 47.72, 46.52, 45.48, 43.8, 42.68, 41.6, 40.24, 39.12, 38.12, 37.0, 35.72, 34.64, 33.72, 32.28, 31.12, 30.08, 29.08, 27.68, 26.56, 25.56, 24.28, 23.16, 22.2, 21.08, 19.88, 18.8, 17.84, 16.56, 15.44, 14.32, 13.32, 12.0, 10.88, 9.96, 7.48, 6.48, 5.4, 4.12, 3.08, 2.08, 1.04}
    pres_qc = 
      {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
    psal = 
      {34.0, 34.0, 34.0, 34.0, 34.0, 33.872, 33.856, 33.848, 33.849, 33.844, 33.839, 33.831, 33.829, 33.826, 33.825, 33.824, 33.822, 33.822, 33.815, 33.807, 33.805, 33.79, 33.783, 33.767, 33.755, 33.75, 33.742, 33.74, 33.735, 33.731, 33.728, 33.723, 33.706, 33.644, 33.593, 33.562, 33.547, 33.518, 33.509, 33.502, 33.478, 33.454, 33.44, 33.441, 33.441, 33.44, 33.439, 33.437, 33.427, 33.414, 33.401, 33.346, 33.335, 33.326, 33.308, 33.245, 33.225, 33.192, 33.121, 33.06, 32.996, 32.94, 32.936, 32.899, 32.879, 32.828, 32.784, 32.773, 32.767, 32.76, 32.756, 32.753, 32.752, 32.751, 32.751, 32.751, 32.749, 32.747, 32.743, 32.723, 32.71, 32.699, 32.696, 32.683, 32.652, 32.648, 32.638, 32.636, 32.631, 32.629, 32.623, 32.618, 32.614, 32.597, 32.594, 32.593, 32.596, 32.589, 32.574, 32.55, 32.555, 33.847, 33.847, 33.847, 33.846, 33.845, 33.846, 33.844, 33.844, 33.842, 33.837, 33.824, 33.815, 33.789, 33.774, 33.768, 33.761, 33.757, 33.753, 33.752, 33.741, 33.7, 33.683, 33.651, 33.652, 33.631, 33.625, 33.618, 33.605, 33.588, 33.572, 33.564, 33.555, 33.552, 33.548, 33.536, 33.512, 33.509, 33.509, 33.503, 33.478, 33.453, 33.44, 33.428, 33.427, 33.404, 33.397, 33.331, 33.269, 33.263, 33.214, 33.141, 33.064, 33.023, 32.962, 32.939, 32.934, 32.932, 32.931, 32.905, 32.867, 32.818, 32.785, 32.774, 32.769, 32.767, 32.764, 32.76, 32.753, 32.741, 32.729, 32.712, 32.695, 32.691, 32.678, 32.645, 32.606, 32.574, 32.558, 32.56, 32.56, 32.56, 32.56, 32.558, 32.559, 32.558, 32.558, 32.556, 32.558, 32.557, 33.855, 33.855, 33.854, 33.849, 33.834, 33.823, 33.82, 33.803, 33.785, 33.775, 33.767, 33.763, 33.761, 33.755, 33.755, 33.755, 33.757, 33.758, 33.757, 33.746, 33.724, 33.706, 33.667, 33.651, 33.634, 33.617, 33.613, 33.608, 33.603, 33.602, 33.598, 33.593, 33.579, 33.555, 33.535, 33.524, 33.505, 33.491, 33.451, 33.431, 33.434, 33.433, 33.423, 33.4, 33.379, 33.338, 33.258, 33.211, 33.164, 33.135, 33.12, 33.112, 33.109, 33.109, 33.109, 33.11, 33.107, 33.045, 32.985, 32.939, 32.938, 32.94, 32.94, 32.89, 32.872, 32.831, 32.784, 32.768, 32.759, 32.753, 32.742, 32.726, 32.713, 32.698, 32.644, 32.592, 32.568, 32.554, 32.551, 32.55, 32.551, 32.548, 32.548, 32.547, 32.546, 32.547, 32.548, 32.545, 32.546, 33.806, 33.803, 33.787, 33.774, 33.758, 33.752, 33.751, 33.75, 33.747, 33.728, 33.711, 33.701, 33.693, 33.681, 33.672, 33.669, 33.667, 33.655, 33.646, 33.633, 33.623, 33.61, 33.6, 33.599, 33.587, 33.583, 33.577, 33.574, 33.57, 33.569, 33.556, 33.547, 33.541, 33.535, 33.529, 33.519, 33.508, 33.501, 33.472, 33.458, 33.444, 33.409, 33.359, 33.289, 33.256, 33.237, 33.196, 33.164, 33.144, 33.131, 33.122, 33.103, 33.075, 33.043, 33.044, 33.017, 33.003, 33.003, 32.981, 32.968, 32.95, 32.915, 32.904, 32.871, 32.846, 32.828, 32.819, 32.812, 32.805, 32.788, 32.782, 32.778, 32.766, 32.753, 32.732, 32.72, 32.679, 32.632, 32.581, 32.559, 32.555, 32.549, 32.549, 32.55, 32.549, 32.549, 32.55, 32.549, 32.549, 32.546, 32.546, 32.546, 32.544}
    psal_qc = 
      {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
    temp = 
      {10.133, 11.679, 12.906, 14.508, 15.446, 9.502, 9.564, 9.614, 9.628, 9.662, 9.695, 9.71, 9.719, 9.725, 9.729, 9.733, 9.739, 9.74, 9.756, 9.765, 9.769, 9.793, 9.796, 9.809, 9.82, 9.822, 9.818, 9.82, 9.824, 9.839, 9.846, 9.854, 9.836, 9.765, 9.713, 9.763, 9.769, 9.837, 9.895, 9.93, 9.999, 10.102, 10.17, 10.186, 10.198, 10.225, 10.255, 10.282, 10.336, 10.39, 10.417, 10.498, 10.501, 10.516, 10.537, 10.558, 10.588, 10.555, 10.414, 10.321, 10.39, 10.312, 10.621, 10.852, 10.951, 10.944, 10.909, 10.908, 10.909, 10.9, 10.892, 10.888, 10.887, 10.886, 10.886, 10.886, 10.888, 10.889, 10.883, 10.876, 10.885, 10.902, 10.915, 10.948, 11.013, 11.025, 11.06, 11.07, 11.082, 11.088, 11.106, 11.126, 11.143, 11.187, 11.196, 11.194, 11.191, 11.212, 11.275, 11.304, 11.287, 9.647, 9.65, 9.653, 9.658, 9.663, 9.666, 9.669, 9.675, 9.685, 9.705, 9.737, 9.761, 9.79, 9.804, 9.811, 9.834, 9.861, 9.893, 9.908, 9.905, 9.84, 9.798, 9.727, 9.73, 9.716, 9.718, 9.729, 9.73, 9.734, 9.755, 9.768, 9.788, 9.793, 9.804, 9.836, 9.904, 9.916, 9.925, 9.942, 10.03, 10.134, 10.23, 10.323, 10.362, 10.425, 10.443, 10.467, 10.446, 10.446, 10.446, 10.317, 10.236, 10.248, 10.257, 10.26, 10.356, 10.632, 10.755, 10.872, 10.914, 10.917, 10.903, 10.898, 10.89, 10.884, 10.881, 10.885, 10.872, 10.868, 10.87, 10.893, 10.935, 10.948, 10.977, 11.069, 11.17, 11.262, 11.312, 11.314, 11.326, 11.332, 11.339, 11.354, 11.358, 11.39, 11.379, 11.399, 11.402, 11.411, 9.623, 9.625, 9.629, 9.647, 9.703, 9.735, 9.744, 9.771, 9.796, 9.806, 9.817, 9.827, 9.833, 9.845, 9.854, 9.862, 9.87, 9.898, 9.912, 9.893, 9.837, 9.797, 9.735, 9.709, 9.699, 9.701, 9.703, 9.703, 9.701, 9.699, 9.697, 9.703, 9.719, 9.767, 9.833, 9.859, 9.921, 9.971, 10.131, 10.315, 10.33, 10.356, 10.405, 10.453, 10.473, 10.475, 10.419, 10.364, 10.305, 10.27, 10.265, 10.258, 10.256, 10.252, 10.252, 10.251, 10.247, 10.216, 10.186, 10.24, 10.24, 10.246, 10.513, 10.729, 10.843, 10.891, 10.897, 10.873, 10.873, 10.861, 10.861, 10.882, 10.906, 10.936, 11.074, 11.206, 11.254, 11.293, 11.308, 11.335, 11.346, 11.369, 11.371, 11.388, 11.408, 11.418, 11.43, 11.454, 11.465, 9.791, 9.794, 9.805, 9.811, 9.817, 9.868, 9.88, 9.898, 9.905, 9.87, 9.816, 9.784, 9.762, 9.744, 9.732, 9.723, 9.721, 9.705, 9.693, 9.689, 9.693, 9.707, 9.721, 9.729, 9.775, 9.789, 9.809, 9.819, 9.835, 9.843, 9.879, 9.903, 9.917, 9.915, 9.919, 9.943, 9.965, 9.989, 10.113, 10.267, 10.368, 10.432, 10.444, 10.424, 10.38, 10.364, 10.32, 10.292, 10.324, 10.352, 10.368, 10.464, 10.448, 10.376, 10.412, 10.84, 10.796, 10.792, 10.808, 10.808, 10.823, 10.889, 10.912, 10.917, 10.908, 10.903, 10.9, 10.897, 10.896, 10.883, 10.876, 10.872, 10.865, 10.86, 10.879, 10.902, 10.999, 11.11, 11.226, 11.293, 11.304, 11.309, 11.318, 11.321, 11.337, 11.342, 11.366, 11.374, 11.406, 11.437, 11.444, 11.461, 11.517}
    temp_qc = 
      {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
    cndc = 
      {3.72344, 3.86723, 3.9826, 4.13482, 4.22476, 3.65783, 3.66195, 3.66572, 3.66709, 3.66968, 3.67219, 3.67275, 3.67334, 3.67356, 3.6738, 3.67401, 3.67433, 3.67438, 3.67513, 3.67512, 3.67525, 3.6759, 3.67543, 3.67498, 3.67475, 3.67439, 3.67318, 3.67311, 3.67293, 3.67383, 3.67412, 3.67431, 3.67094, 3.65833, 3.64855, 3.65002, 3.64905, 3.65236, 3.6567, 3.65915, 3.66303, 3.66999, 3.67475, 3.67626, 3.67731, 3.6796, 3.68218, 3.6844, 3.68828, 3.69187, 3.693, 3.69486, 3.694, 3.69443, 3.6945, 3.69008, 3.69077, 3.68443, 3.66452, 3.64999, 3.64981, 3.63718, 3.66458, 3.68168, 3.68856, 3.68274, 3.67509, 3.67383, 3.67327, 3.67168, 3.6705, 3.66979, 3.66953, 3.66928, 3.66923, 3.66917, 3.66909, 3.66893, 3.66793, 3.66523, 3.66469, 3.66505, 3.66587, 3.66748, 3.67014, 3.67076, 3.67284, 3.67349, 3.674, 3.67429, 3.67526, 3.67651, 3.67759, 3.67975, 3.68021, 3.67988, 3.67987, 3.68101, 3.68509, 3.68521, 3.68415, 3.66857, 3.66883, 3.66907, 3.66939, 3.66972, 3.67006, 3.67011, 3.67061, 3.6713, 3.67261, 3.67423, 3.67551, 3.6756, 3.67536, 3.67538, 3.67675, 3.67879, 3.68126, 3.68248, 3.68106, 3.67104, 3.66548, 3.65582, 3.65614, 3.65275, 3.65229, 3.65254, 3.6513, 3.64995, 3.65023, 3.65057, 3.65143, 3.65154, 3.65209, 3.65376, 3.65754, 3.65829, 3.65903, 3.65993, 3.66544, 3.67239, 3.6798, 3.68705, 3.69045, 3.69386, 3.69477, 3.69034, 3.68221, 3.68158, 3.67665, 3.65765, 3.64265, 3.63962, 3.63433, 3.63226, 3.64036, 3.66498, 3.67592, 3.68383, 3.68374, 3.67901, 3.67437, 3.67274, 3.67146, 3.67067, 3.67002, 3.66992, 3.668, 3.66637, 3.66529, 3.6656, 3.66761, 3.66832, 3.66957, 3.67445, 3.67952, 3.68449, 3.68731, 3.68763, 3.68865, 3.68915, 3.6897, 3.6908, 3.6912, 3.69392, 3.69288, 3.69443, 3.69484, 3.6955, 3.66724, 3.66741, 3.66766, 3.6688, 3.67245, 3.67428, 3.67478, 3.67556, 3.67606, 3.67597, 3.67616, 3.67664, 3.67696, 3.67743, 3.67821, 3.6789, 3.67978, 3.68236, 3.68349, 3.68059, 3.67324, 3.66777, 3.65823, 3.65424, 3.65161, 3.65005, 3.64979, 3.64925, 3.64851, 3.64817, 3.64755, 3.64754, 3.64757, 3.64955, 3.65354, 3.65477, 3.6585, 3.66159, 3.67217, 3.68688, 3.68848, 3.6907, 3.6941, 3.69613, 3.6958, 3.69184, 3.67874, 3.66901, 3.65894, 3.65285, 3.65085, 3.64937, 3.64884, 3.64841, 3.64835, 3.64831, 3.64758, 3.63858, 3.6299, 3.63014, 3.62999, 3.63068, 3.65467, 3.6691, 3.67753, 3.67767, 3.67343, 3.6696, 3.66864, 3.66689, 3.66573, 3.66594, 3.66674, 3.66788, 3.67477, 3.68132, 3.68315, 3.68517, 3.68616, 3.68843, 3.68947, 3.69116, 3.69127, 3.69265, 3.69429, 3.69524, 3.69638, 3.69817, 3.69922, 3.67777, 3.67774, 3.67715, 3.6764, 3.67535, 3.67941, 3.68038, 3.6819, 3.68221, 3.67711, 3.67046, 3.66652, 3.66369, 3.66083, 3.65881, 3.65766, 3.65723, 3.65453, 3.65251, 3.65081, 3.65015, 3.65012, 3.65037, 3.65095, 3.65393, 3.65476, 3.65594, 3.6565, 3.65751, 3.65809, 3.66003, 3.66128, 3.66192, 3.66106, 3.66078, 3.66191, 3.66277, 3.66422, 3.67259, 3.68519, 3.69297, 3.69526, 3.69132, 3.68249, 3.67514, 3.67174, 3.66363, 3.65785, 3.6587, 3.65988, 3.66038, 3.66712, 3.66282, 3.65308, 3.65639, 3.69234, 3.6869, 3.68649, 3.68567, 3.68432, 3.68383, 3.68623, 3.68714, 3.68422, 3.68085, 3.67853, 3.6773, 3.67628, 3.67544, 3.6725, 3.67121, 3.67041, 3.66851, 3.66671, 3.66626, 3.66707, 3.67161, 3.67679, 3.682, 3.68573, 3.68626, 3.68605, 3.68682, 3.68713, 3.68842, 3.68883, 3.69098, 3.69155, 3.69438, 3.69681, 3.69739, 3.69888, 3.70367}
    cndc_qc = 
      {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
    chla = 
      {0.228, 0.228, 0.231, 0.219, 0.216, 0.192, 0.189, 0.189, 0.195, 0.192, 0.192, 0.192, 0.189, 0.192, 0.189, 0.189, 0.192, 0.192, 0.195, 0.192, 0.192, 0.192, 0.189, 0.195, 0.192, 0.192, 0.198, 0.198, 0.195, 0.195, 0.192, 0.195, 0.198, 0.192, 0.198, 0.201, 0.198, 0.195, 0.198, 0.198, 0.201, 0.198, 0.201, 0.201, 0.201, 0.201, 0.198, 0.204, 0.198, 0.201, 0.198, 0.207, 0.207, 0.21, 0.216, 0.219, 0.222, 0.234, 0.243, 0.249, 0.288, 0.339, 0.366, 0.387, 0.408, 0.417, 0.408, 0.432, 0.435, 0.429, 0.42, 0.417, 0.405, 0.417, 0.426, 0.411, 0.438, 0.414, 0.42, 0.426, 0.429, 0.435, 0.426, 0.447, 0.435, 0.429, 0.45, 0.42, 0.432, 0.435, 0.426, 0.417, 0.396, 0.372, 0.351, 0.339, 0.318, 0.294, 0.285, 0.276, 0.276, 0.189, 0.186, 0.192, 0.189, 0.189, 0.195, 0.186, 0.192, 0.189, 0.189, 0.189, 0.189, 0.192, 0.192, 0.192, 0.192, 0.192, 0.195, 0.195, 0.192, 0.201, 0.195, 0.195, 0.195, 0.198, 0.195, 0.192, 0.195, 0.198, 0.195, 0.195, 0.195, 0.195, 0.201, 0.198, 0.198, 0.201, 0.198, 0.201, 0.198, 0.195, 0.195, 0.198, 0.195, 0.201, 0.201, 0.213, 0.21, 0.204, 0.216, 0.222, 0.234, 0.249, 0.261, 0.291, 0.33, 0.351, 0.375, 0.396, 0.396, 0.417, 0.402, 0.411, 0.408, 0.387, 0.384, 0.39, 0.39, 0.411, 0.417, 0.435, 0.456, 0.453, 0.456, 0.423, 0.411, 0.393, 0.366, 0.375, 0.36, 0.357, 0.345, 0.339, 0.312, 0.312, 0.291, 0.288, 0.276, 0.267, 0.192, 0.192, 0.186, 0.189, 0.189, 0.186, 0.192, 0.192, 0.189, 0.189, 0.189, 0.192, 0.192, 0.192, 0.189, 0.192, 0.192, 0.192, 0.189, 0.189, 0.189, 0.192, 0.195, 0.192, 0.192, 0.192, 0.192, 0.192, 0.189, 0.192, 0.195, 0.192, 0.195, 0.192, 0.192, 0.198, 0.198, 0.198, 0.195, 0.198, 0.198, 0.198, 0.201, 0.204, 0.198, 0.204, 0.21, 0.213, 0.222, 0.216, 0.222, 0.225, 0.222, 0.216, 0.219, 0.222, 0.228, 0.246, 0.273, 0.273, 0.27, 0.294, 0.333, 0.354, 0.369, 0.378, 0.411, 0.375, 0.402, 0.39, 0.408, 0.423, 0.462, 0.462, 0.444, 0.423, 0.414, 0.378, 0.375, 0.366, 0.351, 0.324, 0.315, 0.297, 0.288, 0.276, 0.27, 0.255, 0.258, 0.192, 0.186, 0.192, 0.189, 0.186, 0.192, 0.189, 0.189, 0.189, 0.195, 0.192, 0.192, 0.186, 0.189, 0.186, 0.192, 0.192, 0.189, 0.195, 0.192, 0.192, 0.189, 0.192, 0.192, 0.189, 0.192, 0.192, 0.192, 0.189, 0.189, 0.192, 0.195, 0.192, 0.192, 0.195, 0.195, 0.195, 0.192, 0.192, 0.195, 0.192, 0.198, 0.198, 0.201, 0.204, 0.207, 0.213, 0.219, 0.237, 0.231, 0.231, 0.243, 0.249, 0.255, 0.318, 0.333, 0.327, 0.339, 0.339, 0.351, 0.381, 0.39, 0.381, 0.39, 0.381, 0.399, 0.381, 0.396, 0.426, 0.39, 0.396, 0.405, 0.408, 0.426, 0.447, 0.48, 0.474, 0.438, 0.42, 0.411, 0.429, 0.405, 0.387, 0.384, 0.363, 0.327, 0.312, 0.294, 0.288, 0.273, 0.273, 0.261, 0.252}
    chla_qc = 
      {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
    doxy = 
      {281.3286, 271.566, 266.1686, 259.3934, 253.1995, 150.1627, 140.7665, 135.0039, 130.2885, 127.3307, 125.591, 124.3805, 123.7724, 123.3152, 123.0861, 122.9296, 122.929, 123.0763, 123.4629, 123.8468, 124.6823, 125.5296, 126.9756, 128.3544, 129.6549, 130.795, 131.9358, 133.0729, 134.2894, 135.2011, 135.9598, 137.0258, 139.2367, 143.3063, 149.2002, 153.3528, 156.6391, 160.4197, 162.6497, 164.262, 166.7454, 168.2479, 169.4996, 170.7171, 171.8571, 172.3524, 172.6611, 172.8945, 173.3745, 174.0123, 175.1756, 177.6312, 179.3946, 181.0844, 184.5439, 187.4522, 190.5378, 194.613, 200.6862, 205.0068, 211.314, 218.0895, 225.0267, 232.0703, 240.4886, 249.6433, 254.9023, 258.5113, 262.6507, 264.4027, 265.6957, 267.22, 267.7415, 268.1884, 268.5602, 268.9269, 269.0725, 269.2179, 269.5138, 269.6899, 269.9382, 270.261, 270.6453, 270.9841, 271.4468, 271.7552, 272.2398, 272.3525, 272.5074, 272.6175, 272.9359, 272.8293, 272.7203, 272.9521, 272.9895, 273.0543, 273.0366, 272.5531, 272.64, 272.7693, 272.5479, 123.8221, 122.3376, 121.3076, 120.7356, 120.3916, 120.0837, 119.9687, 119.8513, 119.8517, 120.2371, 120.9364, 121.8966, 123.9013, 125.5491, 127.1879, 128.4889, 130.1311, 130.9716, 132.112, 133.7878, 136.6202, 140.0444, 143.0572, 145.6763, 148.0845, 150.4063, 152.2343, 153.8013, 156.2503, 157.8634, 159.5815, 160.8051, 161.6016, 162.7053, 163.7096, 164.7795, 165.8459, 166.4472, 166.9844, 168.3318, 169.3402, 170.0664, 171.2495, 172.0933, 173.2803, 175.4242, 178.5603, 181.8317, 185.5739, 189.9827, 194.6092, 200.562, 206.3492, 212.0908, 216.6283, 222.0206, 227.4092, 231.8155, 239.1746, 245.5246, 251.0385, 256.5952, 260.1976, 262.4871, 264.7747, 265.9868, 266.9025, 267.6644, 268.2062, 268.5243, 269.2481, 270.0543, 270.4398, 271.0056, 271.0267, 271.0656, 271.0107, 271.208, 271.1895, 271.3369, 271.6351, 271.6213, 271.8897, 271.8362, 272.1856, 272.2055, 272.2859, 272.307, 272.378, 122.5643, 121.2323, 120.2047, 119.7924, 120.159, 120.8198, 121.5447, 122.6661, 124.2454, 125.9661, 127.3039, 128.5998, 129.6647, 130.5817, 131.2643, 131.7179, 132.0557, 132.2037, 132.9246, 134.1007, 135.8881, 138.705, 141.6878, 144.8117, 148.8915, 151.1456, 152.6275, 154.3765, 155.6284, 156.3817, 157.33, 158.1277, 159.0542, 160.9176, 162.3231, 163.4398, 165.3792, 166.3908, 167.9314, 169.4915, 170.2451, 171.1617, 172.0176, 173.7314, 175.6612, 178.3756, 183.4135, 187.6454, 191.5726, 195.8681, 198.8553, 200.7639, 202.7442, 203.7994, 204.3995, 205.0752, 206.2106, 209.5646, 214.8305, 219.1166, 221.9368, 224.2956, 228.8346, 233.9008, 242.4692, 248.9811, 254.5714, 258.4826, 261.933, 263.9141, 265.761, 267.1654, 268.1092, 269.0617, 269.5303, 269.7636, 270.0544, 270.856, 270.7017, 271.0114, 271.1573, 271.5409, 271.7172, 271.8687, 271.8679, 272.1658, 272.2362, 272.2021, 272.4237, 129.299, 128.4255, 128.4401, 129.4024, 130.3286, 131.3343, 132.0574, 132.5546, 133.6214, 135.2632, 137.583, 139.4832, 141.1173, 142.7946, 144.2033, 145.6836, 147.3537, 148.5327, 150.2456, 151.5445, 152.8066, 154.152, 155.265, 156.1382, 157.0351, 157.8749, 158.6799, 159.2871, 159.7461, 160.4277, 161.0164, 161.7119, 162.8207, 163.5382, 164.4517, 165.1842, 165.8815, 166.9945, 167.5557, 168.4155, 169.5262, 171.4859, 173.985, 179.0963, 182.8537, 185.7645, 190.1473, 193.3003, 196.767, 199.6111, 201.53, 205.5599, 208.8691, 211.4767, 215.7616, 222.2434, 226.2151, 230.4112, 233.962, 236.575, 240.1998, 244.9499, 248.3363, 251.8326, 256.1145, 258.8111, 260.9589, 262.5682, 264.4087, 265.5687, 266.369, 267.2067, 267.902, 268.2957, 269.0253, 269.5083, 270.2003, 270.0693, 270.5632, 271.0107, 271.1275, 271.3217, 271.8146, 271.8385, 272.0671, 272.2902, 272.3127, 272.3466, 272.4284, 272.6286, 272.7363, 272.6578, 272.4112}
    doxy_qc = 
      {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
    time_gps = 
      {-999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0}
    longitude_gps = 
      {-999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0}
    latitude_gps = 
      {-999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0}
    gps_start_qc = 
      {0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0}
    gps_start_qc_tests = 
      {0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0}
    time_gps_end = 
      {1.6753619999999988E9, 1.6753650000000012E9, 1.6753680000000033E9, 1.6753709999999955E9, 1.6753741200000007E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9}
    latitude_gps_end = 
      {38.3187, 38.3187, 38.3188, 38.3187, 38.3187, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457}
    longitude_gps_end = 
      {-123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693}
    gps_end_qc = 
      {0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0}
    gps_end_qc_tests = 
      {0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0}
    wmo_identifier =   "4801921"
    sensor_doxy = -127
    sensor_ctd = -127
    sensor_fchl = -127
    platform_model =   "Scripps Institution of Oceanography Spray glider"
    platform_serial_number =   "sp028"
    platform_meta = -127
    deployment_time = 
      {1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9}
    deployment_latitude = 
      {38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187}
    deployment_longitude = 
      {-123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713}
}

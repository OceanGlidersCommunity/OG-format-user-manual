netcdf sp041_20191205T1757 {
dimensions:
	N_PARAM = 5 ;
	N_MEASUREMENTS = 25 ;
variables:
	string TRAJECTORY ;
        TRAJECTORY:cf_role = "trajectory_id";
		TRAJECTORY:long_name = "trajectory name";
	string PARAMETER(N_PARAM) ;
		PARAMETER:long_name = "name of parameter computed from glider measurements" ;
		PARAMETER:parameter_vocabulary = "https://vocab.nerc.ac.uk/collection/OG1/current/" ;
	double TIME_GPS(N_MEASUREMENTS) ;
		TIME_GPS:_FillValue = -1. ;
		TIME_GPS:long_name = "time of each GPS location" ;
		TIME_GPS:units = "seconds since 1970-01-01T00:00:00Z" ;
		TIME_GPS:ancillary_variables = "TIME_GPS_QC" ;
      TIME_GPS:calendar = "gregorian" ;
      TIME_GPS:valid_min = 1e9 ;
      TIME_GPS:valid_max = 4e9 ;
	double LATITUDE_GPS(N_MEASUREMENTS) ;
		LATITUDE_GPS:_FillValue = NaN ;
		LATITUDE_GPS:long_name = "latitude of each GPS location" ;
		LATITUDE_GPS:standard_name = "latitude" ;
		LATITUDE_GPS:units = "degrees_north" ;
		LATITUDE_GPS:ancillary_variables = "LATITUDE_GPS_QC" ;
		LATITUDE_GPS:valid_max = "90" ;
		LATITUDE_GPS:valid_min = "-90" ;
	double LONGITUDE_GPS(N_MEASUREMENTS) ;
		LONGITUDE_GPS:_FillValue = NaN ;
		LONGITUDE_GPS:long_name = "longitude of each GPS location" ;
		LONGITUDE_GPS:standard_name = "longitude" ;
		LONGITUDE_GPS:units = "degrees_east" ;
		LONGITUDE_GPS:ancillary_variables = "LONGITUDE_GPS_QC" ;
		LONGITUDE_GPS:valid_max = "180" ;
		LONGITUDE_GPS:valid_min = "-180" ;
	byte PHASE(N_MEASUREMENTS) ;
		PHASE:_FillValue = 0b ;
		PHASE:long_name = "behavior of the glider at sea" ;
		PHASE:ancillary_variables = "PHASE_QC" ;
		PHASE:phase_vocabulary = "url to phase vocab list" ;
		PHASE:phase_calculation_method = "TBD";
		PHASE:phase_calculation_method_vocabulary = "TBD";
		PHASE:phase_calculation_method_doi = "TBD";
	byte PHASE_QC(N_MEASUREMENTS) ;
		PHASE_QC:_FillValue = 0b ;
		PHASE_QC:long_name = "quality flag" ;
	double TIME(N_MEASUREMENTS) ;
		TIME:_FillValue = -1. ;
		TIME:long_name = "time of measurement and GPS location" ;
		TIME:standard_name = "time" ;
		TIME:calendar = "gregorian" ;
		TIME:units = "seconds since 1970-01-01T00:00:00Z" ;
		TIME:valid_min = 1e9 ;
      TIME:valid_max = 4e9 ;
		TIME:interpolation_methodology = "TBD" ;
		TIME:interpolation_methodology_vocabulary = "TBD" ;
		TIME:interpolation_methodology_doi = "TBD" ;
	double LATITUDE(N_MEASUREMENTS) ;
		LATITUDE:_FillValue = -9999.9 ;
		LATITUDE:long_name = "latitude of each measurement and GPS location" ;
		LATITUDE:standard_name = "latitude" ;
		LATITUDE:units = "degrees_north" ;
		LATITUDE:valid_max = "90" ;
		LATITUDE:valid_min = "-90" ;
		LATITUDE:interpolation_methodology = "TBD" ;
		LATITUDE:interpolation_methodology_vocabulary = "TBD" ;
      LATITUDE:interpolation_methodology_doi = "TBD" ;
	double LONGITUDE(N_MEASUREMENTS) ;
		LONGITUDE:_FillValue = -9999.9 ;
		LONGITUDE:long_name = "longitude of each measurements and gps locations" ;
		LONGITUDE:standard_name = "longitude" ;
		LONGITUDE:units = "degrees_east" ;
		LONGITUDE:valid_max = "180" ;
		LONGITUDE:valid_min = "-180" ;
      LONGITUDE:interpolation_methodology = "TBD" ;
      LONGITUDE:interpolation_methodology_vocabulary = "TBD" ;
      LONGITUDE:interpolation_methodology_doi = "TBD" ;
	float PRES(N_MEASUREMENTS) ;
		PRES:_FillValue = -9999.9 ;
		PRES:long_name = "Pressure" ;
		PRES:vocabulary = "http://vocab.nerc.ac.uk/collection/OG1/current/PRES/";
		PRES:standard_name = "sea_water_pressure" ;
		PRES:units = "dbar" ;
		PRES:ancillary_variables = "PRES_QC" ;
		PRES:comment = "Sea water pressure, equals 0 at sea-level" ;
        PRES:sensor = "/CTD";
	byte PRES_QC(N_MEASUREMENTS) ;
		PRES_QC:_FillValue = 0b ;
		PRES_QC:long_name = "quality flag" ;
	float DEPTH(N_MEASUREMENTS) ;
		DEPTH:_FillValue = NaN ;
		DEPTH:long_name = "Depth" ;
		DEPTH:vocabulary = "http://vocab.nerc.ac.uk/collection/OG1/current/DEPTH/";
		DEPTH:standard_name = "depth" ;
		DEPTH:units = "m" ;
		DEPTH:ancillary_variables = "DEPTH_QC" ;
		DEPTH:positive = "down" ;
        DEPTH:sensor = "/CTD";
	byte DEPTH_QC(N_MEASUREMENTS) ;
		DEPTH_QC:_FillValue = 0b ;
		DEPTH_QC:long_name = "quality flag" ;
	float TEMP(N_MEASUREMENTS) ;
		TEMP:_FillValue = -9999.9 ;
		TEMP:long_name = "Sea Water Temperature" ;
		TEMP:vocabulary = "http://vocab.nerc.ac.uk/collection/OG1/current/TEMP/"
		TEMP:standard_name = "sea_water_temperature" ;
		TEMP:units = "Celsius" ;
		TEMP:ancillary_variables = "TEMP_QC" ;
		TEMP:valid_max = 40. ;
		TEMP:valid_min = -5. ;
		TEMP:coverage_content_type = "physicalMeasurement" ;
		TEMP:coordinates = "time lon lat depth" ;
		TEMP:comment = "Sea temperature in-situ ITS-90 scale" ;
        TEMP:sensor = "/CTD";
	byte TEMP_QC(N_MEASUREMENTS) ;
		TEMP_QC:_FillValue = 0b ;
		TEMP_QC:long_name = "quality flag" ;
	float PSAL(N_MEASUREMENTS) ;
		PSAL:_FillValue = NaN ;
		PSAL:long_name = "Sea Water Salinity" ;
		PSAL:vocabulary = "http://vocab.nerc.ac.uk/collection/OG1/current/PSAL/"
		PSAL:standard_name = "sea_water_practical_salinity" ;
		PSAL:units = "1" ;
		PSAL:ancillary_variables = "PSAL_QC" ;
		PSAL:valid_max = 40. ;
		PSAL:valid_min = 0. ;
		PSAL:coverage_content_type = "physicalMeasurement" ;
		PSAL:coordinates = "time lon lat depth" ;
		PSAL:comment = "Practical salinity computed using UNESCO 1983 algorithm" ;
        PSAL:sensor = "/CTD";
	byte PSAL_QC(N_MEASUREMENTS) ;
		PSAL_QC:_FillValue = 0b ;
		PSAL_QC:long_name = "quality flag" ;
	float CHLA(N_MEASUREMENTS) ;
		CHLA:_FillValue = NaN ;
		CHLA:long_name = "Chlorophyll-a concentration" ;
		CHLA:vocabulary = "http://vocab.nerc.ac.uk/collection/OG1/current/CHLA/"
		CHLA:standard_name = "mass_concentration_of_chlorophyll_a_in_sea_water" ;
		CHLA:units = "mg m-3" ;
		CHLA:ancillary_variables = "CHLA_QC" ;
		CHLA:coverage_content_type = "physicalMeasurement" ;
		CHLA:coordinates = "time lon lat depth" ;
		CHLA:comment = "In-situ fluorometer with either manufacturer, laboratory or sample calibration applied" ;
        CHLA:sensor = "/FLUOROMETER_CHLA";
	byte CHLA_QC(N_MEASUREMENTS) ;
		CHLA_QC:_FillValue = 0b ;
		CHLA_QC:long_name = "quality flag" ;
	float DOXY(N_MEASUREMENTS) ;
		DOXY:_FillValue = NaN ;
		DOXY:long_name = "Dissolved oxygen" ;
		DOXY:vocabulary = "http://vocab.nerc.ac.uk/collection/OG1/current/DOXY/"
		DOXY:standard_name = "moles_of_oxygen_per_unit_mass_in_sea_water" ;
		DOXY:units = "micromol kg-1" ;
		DOXY:ancillary_variables = "DOXY_QC" ;
		DOXY:valid_max = 0. ;
		DOXY:valid_min = 500. ;
		DOXY:coverage_content_type = "physicalMeasurement" ;
		DOXY:comment = "Concentration of dissolved oxygen per unit mass of the water column. Oxygen may be expressed in terms of mass, volume or quantity of substance" ;
        DOXY:sensor = "/OPTODE_DOXY";
	byte DOXY_QC(N_MEASUREMENTS) ;
		DOXY_QC:_FillValue = 0b ;
		DOXY_QC:long_name = "quality flag" ;
	double DEPLOYMENT_TIME ;
		DEPLOYMENT_TIME:long_name = "date of deployment" ;
		DEPLOYMENT_TIME:standard_name = "time" ;
		DEPLOYMENT_TIME:calendar = "gregorian" ;
		DEPLOYMENT_TIME:units = "seconds since 1970-01-01T00:00:00Z" ;
		DEPLOYMENT_TIME:axis = "T" ;
	double DEPLOYMENT_LATITUDE ;
		DEPLOYMENT_LATITUDE:long_name = "latitude of deployment" ;
		DEPLOYMENT_LATITUDE:standard_name = "latitude" ;
		DEPLOYMENT_LATITUDE:units = "degrees_north" ;
		DEPLOYMENT_LATITUDE:valid_max = "90" ;
		DEPLOYMENT_LATITUDE:valid_min = "-90" ;
	double DEPLOYMENT_LONGITUDE ;
		DEPLOYMENT_LONGITUDE:long_name = "longitude of deployment" ;
		DEPLOYMENT_LONGITUDE:standard_name = "longitude" ;
		DEPLOYMENT_LONGITUDE:units = "degrees_east" ;
		DEPLOYMENT_LONGITUDE:valid_max = "180" ;
		DEPLOYMENT_LONGITUDE:valid_min = "-180" ;
	string TELECOM_TYPE ;
		TELECOM_TYPE:long_name = "type of telecommunication systems used by the glider" ;
		TELECOM_TYPE:telecom_type_vocabulary = "TBD" ;
	string TRACKING_SYSTEM ;
		TRACKING_SYSTEM:long_name = "type of tracking systems used by the glider" ;
		TRACKING_SYSTEM:tracking_system_vocabulary = "TBD" ;
	string PLATFORM_TYPE ;
		PLATFORM_TYPE:long_name = "type of glider" ;
		PLATFORM_TYPE:platform_type_vocabulary = "https://vocab.nerc.ac.uk/collection/L06/current/";
	string PLATFORM_MODEL ;
		PLATFORM_MODEL:long_name = "model of the glider" ;
		PLATFORM_MODEL:platform_model_vocabulary = "http://vocab.nerc.ac.uk/collection/B76/current/B7600027/";
	string PLATFORM_MAKER ;
		PLATFORM_MAKER:long_name = "Glider manufacturer" ;
		PLATFORM_MAKER:platform_maker_vocabulary = "TBD" ;
	string PLATFORM_SERIAL_NUMBER ;
		PLATFORM_SERIAL_NUMBER:long_name = "glider serial number" ;
	string PLATFORM_CODE ;
		PLATFORM_CODE:long_name = "nickname of the glider" ;
	int PLATFORM_DEPTH_RATING ;
		PLATFORM_DEPTH_RATING:long_name = "Depth limit in meters of the glider for this mission" ;
	string WMO_IDENTIFIER ;
		WMO_IDENTIFIER:long_name = "wmo id" ;
    int INSTRUMENT_CTD ;
        INSTRUMENT_CTD:_FillValue = -2147483647 ;
        INSTRUMENT_CTD:long_name = "Sea-Bird SBE 41CP CTD" ;
  		INSTRUMENT_CTD:type = "CTD" ;
  		INSTRUMENT_CTD:type_vocabulary = "https://vocab.nerc.ac.uk/collection/L05/current/130/" ;
  		INSTRUMENT_CTD:maker = "Sea-Bird Scientific" ;
  		INSTRUMENT_CTD:maker_vocabulary = "https://vocab.nerc.ac.uk/collection/L35/current/MAN0013/" ;
  		INSTRUMENT_CTD:model = "SBE 41CP CTD " ;
  		INSTRUMENT_CTD:model_vocabulary = "https://vocab.nerc.ac.uk/collection/L22/current/TOOL0669/" ;
  		INSTRUMENT_CTD:serial_number = "75" ;
  		INSTRUMENT_CTD:calibration_date = "2019-10-22T00:00:00Z" ;
    int INSTRUMENT_OPTODE_DOXY ;
        INSTRUMENT_OPTODE_DOXY:_FillValue = -2147483647 ;
  		INSTRUMENT_OPTODE_DOXY:long_name = "Sea-Bird SBE 63 dissolved oxygen sensor" ;
  		INSTRUMENT_OPTODE_DOXY:type = "OPTODE_DOXY" ;
  		INSTRUMENT_OPTODE_DOXY:type_vocabulary = "https://vocab.nerc.ac.uk/collection/L05/current/351/" ;
  		INSTRUMENT_OPTODE_DOXY:maker = "Seabird" ;
  		INSTRUMENT_OPTODE_DOXY:maker_vocabulary = "https://vocab.nerc.ac.uk/collection/L35/current/MAN0013/" ;
  		INSTRUMENT_OPTODE_DOXY:model = "Sea-Bird SBE 63 DO" ;
  		INSTRUMENT_OPTODE_DOXY:model_vocabulary = "https://vocab.nerc.ac.uk/collection/L22/current/TOOL0739/" ;
  		INSTRUMENT_OPTODE_DOXY:serial_number = "631776" ;
  		INSTRUMENT_OPTODE_DOXY:calibration_date = "2019-11-22T00:00:00Z" ;
    int INSTRUMENT_FLUOROMETER_CHLA ;     
        INSTRUMENT_FLUOROMETER_CHLA:_FillValue = -2147483647 ;
  		INSTRUMENT_FLUOROMETER_CHLA:long_name = "Seapoint chlorophyll fluorometer" ;
  		INSTRUMENT_FLUOROMETER_CHLA:type = "FLUOROMETER_CHLA" ;
  		INSTRUMENT_FLUOROMETER_CHLA:type_vocabulary = "https://vocab.nerc.ac.uk/collection/L05/current/113/" ;
  		INSTRUMENT_FLUOROMETER_CHLA:maker = "SEAPOINT" ;
  		INSTRUMENT_FLUOROMETER_CHLA:maker_vocabulary = "https://vocab.nerc.ac.uk/collection/L35/current/MAN0177/" ;
  		INSTRUMENT_FLUOROMETER_CHLA:model = "Seapoint SCF" ;
  		INSTRUMENT_FLUOROMETER_CHLA:model_identifier = "http://vocab.nerc.ac.uk/collection/L22/current/TOOL0119/" ;
  		INSTRUMENT_FLUOROMETER_CHLA:serial_number = "S-5012" ;
  		INSTRUMENT_FLUOROMETER_CHLA:calibration_date = "2019-11-22T00:00:00Z" ;

// global attributes:
		:Conventions = "CF-1.8, ACDD-1.3, OG-1.0" ;
		:title = "California Underwater Glider Network - Line 90" ;
		:platform = "sub-surface gliders" ;
		:platform_vocabulary = "https://vocab.nerc.ac.uk/collection/L06/current/27/" ;
		:keywords = "AUVS > Autonomous Underwater Vehicles, Oceans > Ocean Pressure > Water Pressure, Oceans > Ocean Temperature > Water Temperature, Oceans > Salinity/Density > Conductivity, Oceans > Salinity/Density > Density, Oceans > Salinity/Density > Salinity" ;
		:keywords_vocabulary = "GCMD Science Keywords" ;
		:featureType = "trajectory" ;
		:id = "sp041_20191205T1757_R" ;
		:naming_authority = "edu.ucsd.spray" ;
		:history = "readsat - 2020-05-18T19:31:07Z, fixgps3 - 2020-05-18T19:31:07Z, calcvelsat - 2020-05-18T19:31:07Z, calox - 2021-02-26T11:39:46Z, addoxumolkg - 2021-02-26T11:39:46Z" ;
		:comment = "Dataset for demonstration purposes only. Original dataset truncated for the sake of simplicity" ;
		:processing_level = "Automatic quality control" ;
		:standard_name_vocabulary = "CF Standard Name Table v72" ;
		:date_created = "2021-04-10T01:14:44" ;
		:date_modified = "2021-10-06T18:36:50.099674" ;
		:creator_name = "Instrument Development Group" ;
		:creator_email = "idgdata@ucsd.edu" ;
		:creator_url = "http://spraydata.ucsd.edu" ;
		:creator_type = "group" ;
		:creator_institution = "University of California - San Diego; Scripps Institution of Oceanography" ;
		:institution = "Scripps Institution of Oceanography" ;
		:project = "California Underwater Glider Network" ;
		:publisher_name = "Instrument Development Group" ;
		:publisher_email = "idgdata@ucsd.edu" ;
		:publisher_url = "https://spraydata.ucsd.edu" ;
		:publisher_type = "group" ;
		:publisher_institution = "University of California - San Diego; Scripps Institution of Oceanography" ;
		:geospatial_bounds = "POLYGON ((-119.82769 32.50146, -119.821205 32.50548, -119.80175 32.51754, -119.82769 32.50146))" ;
		:geospatial_bounds_crs = "EPSG:4326" ;
		:geospatial_bounds_vertical_crs = "EPSG:5831" ;
		:geospatial_lat_min = 32.50146 ;
		:geospatial_lat_max = 32.51754 ;
		:geospatial_lon_min = -119.82769 ;
		:geospatial_lon_max = -119.80175 ;
		:geospatial_vertical_min = 1.54 ;
		:geospatial_vertical_max = 24.59 ;
		:geospatial_vertical_positive = "down" ;
		:geospatial_vertical_units = "m" ;
		:time_coverage_start = "2019-12-05T17:57Z" ;
		:time_coverage_end = "2019-12-05T18:05Z" ;
		:program = "GOMO, IOOS" ;
		:network = "California Underwater Glider Network" ;
		:project = "California Underwater Glider Network" ;
		:contributor_name = "Daniel Rudnick,Guilherme Castelao" ;
		:contributor_role = "Principal Investigator, Data Curator" ;
		:product_version = "v3" ;
		:instrument = "Sea-Bird 41CP" ;
		:metadata_link = "http://spraydata.ucsd.edu" ;
		:ctd_make_model = "Sea-Bird 41CP" ;
		:doi = "10.21238/S8SPRAY1618" ;
		:xglider_type = "trajectoryObs" ;
		:trajectory = "sp041_20191205T1757" ;
		:wmoid = "4801948" ;
		:internal_mission_identifier = "19C04101" ;
		:site = "CUGN line 90" ;
		:site_vocabulary = "TBD" ;
		:network = "California Underwater Glider Network" ;
		:contributor_email = "drudnick@ucsd.edu,castelao@ucsd.edu" ;
		:contributor_id = "0000-0002-2624-7074,0000-0002-6765-0708" ;
		:contributor_role_vocabulary = "https://orcid.org/" ;
		:contributor_role = "Principal Investigator, Data Curator" ;
		:agency = "Scripps Institution of Oceanography" ;
		:agency_role = "SDNPR004" ;
		:agency_role_vocabulary = "http://vocab.nerc.ac.uk/collection/C86/" ;
		:agency_id = "1390" ;
		:agency_id_vocabulary = "EDMO" ;
		:data_url = "https://spraydata.ucsd.edu/projects/CUGN/" ;
		:rtqc_method = "Spray - CoTeDe" ;
		:rtqc_method_doi = "10.21105/joss.02063" ;
		:web_link = "https://spraydata.ucsd.edu/projects/CUGN/" ;
		:mission = "19C04101" ;
data:

 TRAJECTORY = "sp041_20191205T1757" ;

 PARAMETER = "PRES", "TEMP", "PSAL", "CHLA", "DOXY" ;

 TIME_GPS = 1576507260, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, 1576517403 ;

 LATITUDE_GPS = 32.51754, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, 32.50146 ;

 LONGITUDE_GPS = -119.80175, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, -119.82769 ;

 PHASE = _, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, _ ;

 PHASE_QC = _, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, _ ;

 TIME = 1576507260, 1576516817, 1576516825, 1576516833, 1576516841, 
    1576516849, 1576516857, 1576516865, 1576516873, 1576516881, 1576516889, 
    1576516897, 1576516905, 1576516913, 1576516921, 1576516929, 1576516937, 
    1576516945, 1576516953, 1576516961, 1576516969, 1576516977, 1576516985, 
    1576516993, 1576517403 ;

 LATITUDE = 32.51754, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, 32.50146 ;

 LONGITUDE = -119.80175, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, -119.82769 ;

 PRES = _, 24.76, 23.68, 22.76, 21.72, 20.72, 19.68, 18.64, 17.48, 16.6, 
    15.52, 14.6, 13.44, 12.44, 11.4, 10.2, 8.44, 7.44, 6.28, 5.32, 4.36, 3.4, 
    2.32, 1.56, _ ;

 PRES_QC = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _ ;

 DEPTH = _, 24.5849769627501, 23.5126728256206, 22.5992241312562, 
    21.5666250478649, 20.5737364026879, 19.5411271039573, 18.5085125971717, 
    17.3567441183672, 16.4829843983173, 15.4106378268966, 14.4971529837432, 
    13.3453619368607, 12.3524334192887, 11.3197826520277, 10.1282560628289, 
    8.38067118597407, 7.38771858618288, 6.23588753584426, 5.28264314410755, 
    4.32939431287006, 3.37614104200687, 2.30372580539014, 1.5490598630261, _ ;

 TEMP = _, 15.505, 15.506, 15.505, 15.505, 15.506, 15.505, 15.505, 15.505, 
    15.504, 15.506, 15.504, 15.505, 15.508, 15.507, 15.509, 15.509, 15.51, 
    15.51, 15.511, 15.51, 15.511, 15.512, 15.512, _ ;

 TEMP_QC = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _ ;

 PSAL = _, 33.561, 33.561, 33.561, 33.561, 33.562, 33.561, 33.561, 33.561, 
    33.562, 33.561, 33.561, 33.561, 33.561, 33.561, 33.561, 33.561, 33.561, 
    33.56, 33.561, 33.56, 33.56, 33.559, 33.56, _ ;

 PSAL_QC = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _ ;

 CHLA = _, 0.861, 0.909, 0.873, 0.867, 0.834, 0.864, 0.882, 0.855, 0.93, 
    0.819, 0.786, 0.807, 0.783, 0.741, 0.744, 0.609, 0.555, 0.573, 0.498, 
    0.471, 0.453, 0.444, 0.414, _ ;

 CHLA_QC = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _ ;

 DOXY = _, 240.699500381006, 240.728111146589, 240.75690836507, 
    240.710612669174, 240.922144300944, 240.655413148225, 240.720151525978, 
    240.635340339479, 240.700230807224, 240.76636985969, 240.831706998232, 
    240.7111499353, 240.664998530651, 240.915858055632, 240.904784287258, 
    241.074164770971, 240.990908679491, 241.093556991221, 241.119569863555, 
    241.297597492548, 241.067163480339, 241.244566377113, 241.199209516033, _ ;

 DOXY_QC = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
    _, _, _ ;

 DEPLOYMENT_TIME = 1575570735.0 ;

 DEPLOYMENT_LATITUDE = 32.9018 ;

 DEPLOYMENT_LONGITUDE = -117.29972500000001 ;

 TELECOM_TYPE = "Iridium" ;

 TRACKING_SYSTEM = "GPS, ARGOS" ;

 PLATFORM_TYPE = "Spray" ;

 PLATFORM_MODEL = "Spray" ;

 PLATFORM_MAKER = "Scripps Institution of Oceanography" ;

 PLATFORM_SERIAL_NUMBER = "0041" ;

 PLATFORM_CODE = "sp041" ;

 PLATFORM_DEPTH_RATING = 1000 ;

 WMO_IDENTIFIER = "4801948" ;

 INSTRUMENT_CTD = _ ;

 INSTRUMENT_OPTODE_DOXY = _ ;

 INSTRUMENT_FLUOROMETER_CHLA = _ ;
}

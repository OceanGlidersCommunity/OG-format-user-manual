netcdf file:/Users/sevadjian/projects/spraydata-dev/erddap_stuff/erddap_data/ocean_gliders/sp028_20230202T1637_R.nc {
  dimensions:
    n_measurements = UNLIMITED;   // (1493 currently)
  variables:
    String trajectory;
      :cf_role = "trajectory_id";
      :comment = "A trajectory is one deployment of a glider. The format is platform_id-YYYYMMDDThhmm. Where the time is the start of the first dive of the trajectory.";
      :long_name = "Trajectory Name";

    int profile_index(n_measurements=1493);
      :ioos_category = "Identifier";
      :long_name = "Profile Number";
      :valid_max = 2147483647; // int
      :valid_min = 1; // int
      :comment = "Sequential profile number within the trajectory, extended for use along the \'obs\' dimension\'. Use this variable for indexing or shaping the data. The first profile has a value of 1 and is incremented for each successive profile contained in the trajectory.";
      :_FillValue = -999; // int
      :_ChunkSizes = 1024U; // uint

    double time_profile(n_measurements=1493);
      :_CoordinateAxisType = "Time";
      :long_name = "Profile Time";
      :axis = "T";
      :calendar = "gregorian";
      :comment = "An estimate of the time of the mid-point of each profile. time_profile = time_gps + 0.75 * (time_gps_end - time_gps);";
      :ioos_category = "Time";
      :observation_type = "calculated";
      :platform = "platform_meta";
      :standard_name = "time";
      :time_origin = "01-JAN-1970 00:00:00";
      :units = "seconds since 1970-01-01T00:00:00Z";
      :ancillary_variables = "time_profile_qc";
      :_ChunkSizes = 512U; // uint

    int time_profile_qc(n_measurements=1493);
      :_FillValue = -127; // int
      :long_name = "Profile Time Quality Flag";
      :standard_name = "aggregate_quality_flag";
      :valid_max = 9; // int
      :valid_min = 0; // int
      :flag_values = 1, 2, 3, 4, 9; // int
      :flag_meanings = "good not_evaluated questionable bad missing";
      :comment = "1=Good/Pass, 2=Not Evaluated, 3=Questionable, Suspect or of High Interest, 4=Fail/Bad, 9=Missing Data. See the references for more details on the flag meanings.";
      :references = "Paris. Intergovernmental Oceanographic Commission of UNESCO, 2013. Ocean Data Standards, Vol.3:Recommendation for a Quality Flag Scheme for the Exchange of Oceanographic and Marine    Meteorological Data. (IOC Manuals and Guides, 54, Vol. 3.) 12 pp. (English.)(IOC/2013/MG/54-3) https://repository.oceanbestpractices.org/bitstream/handle/11329/413/MG54_3.doc";
      :_ChunkSizes = 747U; // uint

    double latitude_profile(n_measurements=1493);
      :_FillValue = -999.0; // double
      :_CoordinateAxisType = "Lat";
      :long_name = "Profile Latitude, Mid-Point";
      :axis = "Y";
      :colorBarMaximum = 90.0; // double
      :colorBarMinimum = -90.0; // double
      :comment = "An estimate of the latitude at the mid-point of each profile. latitude_profile = latitude_gps + 0.75 * (latitude_gps_end - latitude_gps);";
      :ioos_category = "Location";
      :observation_type = "calculated";
      :platform = "platform_meta";
      :standard_name = "latitude";
      :units = "degrees_north";
      :valid_max = 90.0; // double
      :valid_min = -90.0; // double
      :ancillary_variables = "latitude_profile_qc";
      :_ChunkSizes = 498U; // uint

    int latitude_profile_qc(n_measurements=1493);
      :_FillValue = -127; // int
      :long_name = "Profile Latitude Mid-Point Quality Flag";
      :standard_name = "aggregate_quality_flag";
      :valid_max = 9; // int
      :valid_min = 0; // int
      :flag_values = 1, 2, 3, 4, 9; // int
      :flag_meanings = "good not_evaluated questionable bad missing";
      :comment = "1=Good/Pass, 2=Not Evaluated, 3=Questionable, Suspect or of High Interest, 4=Fail/Bad, 9=Missing Data. See the references for more details on the flag meanings.";
      :references = "Paris. Intergovernmental Oceanographic Commission of UNESCO, 2013. Ocean Data Standards, Vol.3:Recommendation for a Quality Flag Scheme for the Exchange of Oceanographic and Marine    Meteorological Data. (IOC Manuals and Guides, 54, Vol. 3.) 12 pp. (English.)(IOC/2013/MG/54-3) https://repository.oceanbestpractices.org/bitstream/handle/11329/413/MG54_3.doc";
      :_ChunkSizes = 747U; // uint

    double latitude_uv(n_measurements=1493);
      :_FillValue = -999.0; // double
      :long_name = "Latitude of Underwater Segment Mid-Point Estimate";
      :axis = "Y";
      :colorBarMaximum = 90.0; // double
      :colorBarMinimum = -90.0; // double
      :comment = "This latitude variable is provided specifically for use with the depth-averaged current variables u and v. The value is an estimate of the glider location at the midpoint of the underwater segment. It differs from the latitude variable which is the estimate of the mid-point of the profile which is at 3/4 of the underwater segment. The value is interpolated to provide an estimate of the mid-point of the entire underwater segment, which may consist of 1 or more dives. Calculated using surface GPS positions at the start and end of the dive. Where, latitude_uv = latitude_gps + 0.5 * (latitude_gps_end - latitude_gps);";
      :ioos_category = "Location";
      :observation_type = "calculated";
      :platform = "platform_meta";
      :standard_name = "latitude";
      :units = "degrees_north";
      :valid_max = 90.0; // double
      :valid_min = -90.0; // double
      :ancillary_variables = "latitude_uv_qc";
      :_ChunkSizes = 498U; // uint

    int latitude_uv_qc(n_measurements=1493);
      :_FillValue = -127; // int
      :long_name = "Latitude of Underwater Segment Mid-Point Estimate Quality Flag";
      :valid_max = 9; // int
      :valid_min = 1; // int
      :flag_values = 1, 2, 3, 4, 9; // int
      :flag_meanings = "good not_evaluated questionable bad missing";
      :comment = "1=Good/Pass, 2=Not Evaluated, 3=Questionable, Suspect or of High Interest, 4=Fail/Bad, 9=Missing Data. See the references for more details on the flag meanings.";
      :references = "Paris. Intergovernmental Oceanographic Commission of UNESCO, 2013. Ocean Data Standards, Vol.3:Recommendation for a Quality Flag Scheme for the Exchange of Oceanographic and Marine    Meteorological Data. (IOC Manuals and Guides, 54, Vol. 3.) 12 pp. (English.)(IOC/2013/MG/54-3) https://repository.oceanbestpractices.org/bitstream/handle/11329/413/MG54_3.doc";
      :_ChunkSizes = 747U; // uint

    double longitude_profile(n_measurements=1493);
      :_FillValue = -999.0; // double
      :long_name = "Profile Mid-Point Longitude";
      :axis = "X";
      :comment = "An estimate of the longitude at the mid-point of each profile. longitude_profile = longitude_gps + 0.75 * (longitude_gps_end - longitude_gps);";
      :ioos_category = "Location";
      :observation_type = "calculated";
      :platform = "platform_meta";
      :standard_name = "longitude";
      :units = "degrees_east";
      :valid_max = 180.0; // double
      :valid_min = -180.0; // double
      :ancillary_variables = "longitude_profile_qc";
      :_ChunkSizes = 498U; // uint

    int longitude_profile_qc(n_measurements=1493);
      :_FillValue = -127; // int
      :long_name = "Profile Longitude Quality Flag";
      :standard_name = "aggregate_quality_flag";
      :valid_max = 9; // int
      :valid_min = 1; // int
      :flag_values = 1, 2, 3, 4, 9; // int
      :flag_meanings = "good not_evaluated questionable bad missing";
      :comment = "1=Good/Pass, 2=Not Evaluated, 3=Questionable, Suspect or of High Interest, 4=Fail/Bad, 9=Missing Data. See the references for more details on the flag meanings.";
      :references = "Paris. Intergovernmental Oceanographic Commission of UNESCO, 2013. Ocean Data Standards, Vol.3:Recommendation for a Quality Flag Scheme for the Exchange of Oceanographic and Marine    Meteorological Data. (IOC Manuals and Guides, 54, Vol. 3.) 12 pp. (English.)(IOC/2013/MG/54-3) https://repository.oceanbestpractices.org/bitstream/handle/11329/413/MG54_3.doc";
      :_ChunkSizes = 747U; // uint

    double longitude_uv(n_measurements=1493);
      :_FillValue = -999.0; // double
      :long_name = "Longitude of Underwater Segment (Mid-Point Estimate)";
      :axis = "X";
      :comment = "This longitude variable is provided specifically for use with the depth-averaged current variables u and v. The value is an estimate of the glider location at the midpoint of the underwater segment. It differs from the longitude_profile variable which is the estimate of the mid-point of the profile which is at 3/4 of the underwater segment. The value is interpolated to provide an estimate of the mid-point of the entire underwater segment, which may consist of 1 or more dives. Calculated using surface GPS positions at the starta nd end of the dive. Where, longitude_uv = longitude_gps + 0.5 * (longitude_gps_end - longitude_gps);";
      :ioos_category = "Location";
      :observation_type = "calculated";
      :platform = "platform_meta";
      :standard_name = "longitude";
      :units = "degrees_east";
      :valid_max = 180.0; // double
      :valid_min = -180.0; // double
      :ancillary_variables = "longitude_uv_qc";
      :_ChunkSizes = 498U; // uint

    int longitude_uv_qc(n_measurements=1493);
      :_FillValue = -127; // int
      :long_name = "Longitude of Underwater Segment (Mid-Point Estimate) Quality Flag";
      :valid_max = 9; // int
      :valid_min = 1; // int
      :flag_values = 1, 2, 3, 4, 9; // int
      :flag_meanings = "good not_evaluated questionable bad missing";
      :comment = "1=Good/Pass, 2=Not Evaluated, 3=Questionable, Suspect or of High Interest, 4=Fail/Bad, 9=Missing Data. See the references for more details on the flag meanings.";
      :references = "Paris. Intergovernmental Oceanographic Commission of UNESCO, 2013. Ocean Data Standards, Vol.3:Recommendation for a Quality Flag Scheme for the Exchange of Oceanographic and Marine    Meteorological Data. (IOC Manuals and Guides, 54, Vol. 3.) 12 pp. (English.)(IOC/2013/MG/54-3) https://repository.oceanbestpractices.org/bitstream/handle/11329/413/MG54_3.doc";
      :_ChunkSizes = 747U; // uint

    double time_uv(n_measurements=1493);
      :_FillValue = -999.0; // double
      :long_name = "Time Estimate for Underwater Segment";
      :axis = "T";
      :comment = "This time variable is provided for use with the depth-averaged current variables u and v. The value is an estimate of the glider location at the midpoint of the underwater segment. The value is interpolated to provide an estimate of the mid-point of the entire underwater segment, which may consist of 1 or more dives. Calculated using surface GPS times at the start and end of the dive. Where, time_uv = time_gps + 0.5 * (time_gps_end - time_gps);";
      :ioos_category = "Time";
      :observation_type = "calculated";
      :platform = "platform_meta";
      :standard_name = "time";
      :units = "seconds since 1970-01-01T00:00:00Z";
      :time_origin = "01-JAN-1970 00:00:00";
      :ancillary_variables = "time_uv_qc";
      :_ChunkSizes = 498U; // uint

    int time_uv_qc(n_measurements=1493);
      :_FillValue = -127; // int
      :coverage_content_type = "qualityInformation";
      :long_name = "Time Estimate for Underwater Segment Quality Flag";
      :valid_max = 9; // int
      :valid_min = 1; // int
      :flag_values = 1, 2, 3, 4, 9; // int
      :flag_meanings = "good not_evaluated questionable bad missing";
      :comment = "1=Good/Pass, 2=Not Evaluated, 3=Questionable, Suspect or of High Interest, 4=Fail/Bad, 9=Missing Data. See the references for more details on the flag meanings.";
      :references = "Paris. Intergovernmental Oceanographic Commission of UNESCO, 2013. Ocean Data Standards, Vol.3:Recommendation for a Quality Flag Scheme for the Exchange of Oceanographic and Marine    Meteorological Data. (IOC Manuals and Guides, 54, Vol. 3.) 12 pp. (English.)(IOC/2013/MG/54-3) https://repository.oceanbestpractices.org/bitstream/handle/11329/413/MG54_3.doc";
      :_ChunkSizes = 747U; // uint

    double time(n_measurements=1493);
      :_FillValue = -999.0; // double
      :_CoordinateAxisType = "Time";
      :long_name = "Time of Each Observation";
      :axis = "T";
      :calendar = "gregorian";
      :comment = "Time stamp at each point in the underwater profile during a dive. This time stamp corresponds to the acquisition of the sensor data.";
      :ioos_category = "Time";
      :observation_type = "measured";
      :platform = "platform_meta";
      :standard_name = "time";
      :time_origin = "01-JAN-1970 00:00:00";
      :units = "seconds since 1970-01-01T00:00:00Z";
      :_ChunkSizes = 498U; // uint

    int time_qc(n_measurements=1493);
      :_FillValue = -127; // int
      :comment = "Subsurface time values are more accurate than subsurface latitude and longitude. Subsurface positions are best estimates with lower accuracy. See the corresponding position variable metadata for more details. 1=Good/Pass, 2=Not Evaluated, 3=Questionable, Suspect or of High Interest, 4=Fail/Bad, 9=Missing Data. See the references for more details on the flag meanings.";
      :coverage_content_type = "qualityInformation";
      :flag_values = 1, 2, 3, 4, 9; // int
      :flag_meanings = "good not_evaluated questionable bad missing";
      :long_name = "Quality Flag for the Time of Each Observation";
      :standard_name = "aggregate_quality_flag";
      :references = "Paris. Intergovernmental Oceanographic Commission of UNESCO, 2013. Ocean Data Standards, Vol.3:Recommendation for a Quality Flag Scheme for the Exchange of Oceanographic and Marine    Meteorological Data. (IOC Manuals and Guides, 54, Vol. 3.) 12 pp. (English.)(IOC/2013/MG/54-3) https://repository.oceanbestpractices.org/bitstream/handle/11329/413/MG54_3.doc";
      :valid_max = 9; // int
      :valid_min = 0; // int
      :_ChunkSizes = 747U; // uint

    double wcur_x(n_measurements=1493);
      :_FillValue = -999.0; // double
      :ancillary_variables = "wcur_qc wcur_qc_tests";
      :colorBarMaximum = 0.5; // double
      :colorBarMinimum = 0.5; // double
      :comment = "The depth-averaged current is an estimate of the net current measured while the glider is underwater. The value is calculated over the entire underwater segment. The latitude_uv, longitude_uv and time_uv variables provide the location and time for this variable. Additional velocity data are available from the acoustic doppler current profiler (ADCP). Please contact us at idgdata@ucsd.edu if you are interested in the ADCP data.";
      :coordinates = "time_uv longitude_uv latitude_uv";
      :coverage_content_type = "physicalMeasurement";
      :ioos_category = "Location";
      :long_name = "U, Depth-Averaged Eastward Sea Water Velocity";
      :observation_type = "calculated";
      :platform = "platform_meta";
      :standard_name = "eastward_sea_water_velocity";
      :units = "m s-1";
      :valid_max = 10.0; // double
      :valid_min = -10.0; // double
      :vocabulary = "https://vocab.nerc.ac.uk/collection/OG1/current";
      :_ChunkSizes = 498U; // uint

    double wcur_y(n_measurements=1493);
      :_FillValue = -999.0; // double
      :ancillary_variables = "wcur_qc wcur_qc_tests";
      :colorBarMaximum = 0.5; // double
      :colorBarMinimum = 0.5; // double
      :comment = "The depth-averaged current is an estimate of the net current measured while the glider is underwater. The value is calculated over the entire underwater segment. The latitude_uv, longitude_uv and time_uv variables provide the location and time for this variable. Additional velocity data are available from the acoustic doppler current profiler (ADCP). Please contact us at idgdata@ucsd.edu if you are interested in the ADCP data.";
      :coordinates = "time_uv longitude_uv latitude_uv";
      :coverage_content_type = "physicalMeasurement";
      :ioos_category = "Location";
      :long_name = "V, Depth-Averaged Northward Sea Water Velocity";
      :observation_type = "calculated";
      :platform = "platform_meta";
      :standard_name = "northward_sea_water_velocity";
      :units = "m s-1";
      :valid_max = 10.0; // double
      :valid_min = -10.0; // double
      :vocabulary = "https://vocab.nerc.ac.uk/collection/OG1/current";
      :_ChunkSizes = 498U; // uint

    int wcur_qc(n_measurements=1493);
      :_FillValue = -127; // int
      :comment = "The depth averaged velocity calculation is dependent on the glider position at the start and end of each dive. These flags are derived from the GPS flags for the dive. 1=Good/Pass, 2=Not Evaluated, 3=Questionable, Suspect or of High Interest, 4=Fail/Bad, 9=Missing Data. See the references for more details on the flag meanings.";
      :coverage_content_type = "qualityInformation";
      :flag_values = 1, 2, 3, 4, 9; // int
      :flag_meanings = "good not_evaluated questionable bad missing";
      :long_name = "Depth-Averaged Sea Water Velocity Quality Flag";
      :standard_name = "aggregate_quality_flag";
      :valid_max = 9; // int
      :valid_min = 1; // int
      :_ChunkSizes = 747U; // uint

    int wcur_qc_tests(n_measurements=1493);
      :_FillValue = -127; // int
      :coverage_content_type = "qualityInformation";
      :long_name = "Depth-Averaged Eastward Sea Water Velocity Quality Flag";
      :valid_max = 99; // int
      :valid_min = 0; // int
      :flag_values = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 99; // int
      :flag_meanings = "gps_good gps_day_problem gps_repeat gps_backward gps_too_fast_on_surface gps_too_soon gps_too_far gps_bad_hdop gps_bad_status gps_no_surfacing gps_manual gps_no_dive";
      :standard_name = "quality_flag";
      :comment = "The depth averaged velocity calculation on the glider position at the start and end of each dive. These flags are derived from the GPS flags for the dive. gps_good=0 gps_day_problem=1 gps_repeat=2 gps_backward=3 gps_too_fast_on_surface=4 gps_too_soon=5 gps_too_far=6 gps_bad_hdop=7 gps_bad_status=8 gps_no_surfacing=9 gps_manual=10 gps_no_dive=99";
      :_ChunkSizes = 747U; // uint

    double depth(n_measurements=1493);
      :_FillValue = -999.0; // double
      :_CoordinateAxisType = "Height";
      :_CoordinateZisPositive = "down";
      :ancillary_variables = "depth_qc";
      :axis = "Z";
      :colorBarMaximum = 2000.0; // double
      :colorBarMinimum = 0.0; // double
      :colorBarPalette = "OceanDepth";
      :ioos_category = "Location";
      :long_name = "Depth";
      :observation_type = "calculated";
      :platform = "platform_meta";
      :positive = "down";
      :reference_datum = "sea-surface";
      :sensor = "sensor_ctd";
      :standard_name = "depth";
      :units = "m";
      :valid_max = 2000.0; // double
      :valid_min = 0.0; // double
      :vocabulary = "https://vocab.nerc.ac.uk/collection/OG1/current";
      :comment = "Depth values are calculated from pressure. A Spray glider profiles on the ascent, collecting sensor data beginning in deeper water and ending at the surface.";
      :_ChunkSizes = 498U; // uint

    int depth_qc(n_measurements=1493);
      :_FillValue = -127; // int
      :comment = "1=Good/Pass, 2=Not Evaluated, 3=Questionable, Suspect or of High Interest, 4=Fail/Bad, 9=Missing Data. See the references for more details on the flag meanings.";
      :coverage_content_type = "qualityInformation";
      :long_name = "Depth Quality Flag";
      :standard_name = "aggregate_quality_flag";
      :flag_values = 1, 2, 3, 4, 9; // int
      :flag_meanings = "good not_evaluated questionable bad missing";
      :references = "Paris. Intergovernmental Oceanographic Commission of UNESCO, 2013. Ocean Data Standards, Vol.3:Recommendation for a Quality Flag Scheme for the Exchange of Oceanographic and Marine    Meteorological Data. (IOC Manuals and Guides, 54, Vol. 3.) 12 pp. (English.)(IOC/2013/MG/54-3) https://repository.oceanbestpractices.org/bitstream/handle/11329/413/MG54_3.doc";
      :valid_max = 9; // int
      :valid_min = 0; // int
      :_ChunkSizes = 747U; // uint

    double latitude(n_measurements=1493);
      :_FillValue = -999.0; // double
      :long_name = "Estimated Subsurface Latitude";
      :colorBarMaximum = 90.0; // double
      :colorBarMinimum = -90.0; // double
      :comment = "Estimated position of the glider underwater during a dive. Use the GPS position variables for accurate positions at the surface. Use caution with these estimated subsurface position values, the deviation from actual position may be several hundreds of meters! Estimations are a dead reckoning using the GPS positions at the start and end of the dive, and the gliders estimated velocity. The calculation methods are described in: \'Rudnick, D. L., Sherman, J. T., & Wu, A. P. (2018). Depth-average velocity from Spray underwater gliders. Journal of Atmospheric and Oceanic Technology, (2018), 35, 1665-1673; doi: https://doi.org/10.1175/JTECH-D-17-0200.1\'. The accuracy attribute reflects an accuracy of approximately +/-800m (0.007 &deg;)";
      :ioos_category = "Location";
      :observation_type = "calculated";
      :platform = "platform_meta";
      :standard_name = "latitude";
      :units = "degrees_north";
      :valid_max = 90.0; // double
      :valid_min = -90.0; // double
      :references = "Rudnick, D. L., Sherman, J. T., & Wu, A. P. (2018). Depth-average velocity from Spray underwater gliders. Journal of Atmospheric and Oceanic Technology, (2018), 35, 1665-1673; doi: https://doi.org/10.1175/JTECH-D-17-0200.1";
      :accuracy = 0.007; // double
      :_ChunkSizes = 498U; // uint

    int latitude_qc(n_measurements=1493);
      :_FillValue = -127; // int
      :coverage_content_type = "qualityInformation";
      :long_name = "Quality Flag for the Estimated Subsurface Latitude";
      :short_name = "Quality Flag for Subsurface Latitude";
      :standard_name = "aggregate_quality_flag";
      :valid_max = 9; // int
      :valid_min = 0; // int
      :flag_values = 1, 2, 3, 4, 9; // int
      :flag_meanings = "good not_evaluated questionable bad missing";
      :comment = "Use caution - these are estimated subsurface position values, the deviation from actual position may be several hundreds of meters! These are estimations and are a dead reckoning using the GPS positions at dive start and end, and the gliders estimated velocity. The calculation methods are described in Rudnick, D. L., Sherman, J. T., & Wu, A. P. (2018). Depth-average velocity from Spray underwater gliders. Journal of Atmospheric and Oceanic Technology, (2018), 35, 1665-1673; doi: https://doi.org/10.1175/JTECH-D-17-0200.1. The accuracy attribute reflects an accuracy of approximately +/-800m (0.09 &deg; Lon) 1=Good/Pass, 2=Not Evaluated, 3=Questionable, Suspect or of High Interest, 4=Fail/Bad, 9=Missing Data. See the references for more details on the flag meanings.";
      :references = "Paris. Intergovernmental Oceanographic Commission of UNESCO, 2013. Ocean Data Standards, Vol.3:Recommendation for a Quality Flag Scheme for the Exchange of Oceanographic and Marine    Meteorological Data. (IOC Manuals and Guides, 54, Vol. 3.) 12 pp. (English.)(IOC/2013/MG/54-3) https://repository.oceanbestpractices.org/bitstream/handle/11329/413/MG54_3.doc";
      :_ChunkSizes = 747U; // uint

    double longitude(n_measurements=1493);
      :_FillValue = -999.0; // double
      :axis = "X";
      :colorBarMaximum = 180.0; // double
      :colorBarMinimum = -180.0; // double
      :comment = "Use caution - these are estimated positions of the glider underwater during a dive. Use the GPS position variables for accurate positions at the surface. Use caution with these estimated subsurface position values, the deviation from actual position may be several hundreds of meters! These estimations are a dead reckoning using the GPS positions at dive start and end, and the gliders estimated velocity. The calculation methods are described in: \'Rudnick, D. L., Sherman, J. T., & Wu, A. P. (2018). Depth-average velocity from Spray underwater gliders. Journal of Atmospheric and Oceanic Technology, (2018), 35, 1665-1673; doi: https://doi.org/10.1175/JTECH-D-17-0200.1\'. The accuracy attribute reflects an accuracy of approximately +/-800m (0.09 &deg; Lon)";
      :ioos_category = "Location";
      :long_name = "Estimated Subsurface Longitude";
      :observation_type = "calculated";
      :platform = "platform_meta";
      :standard_name = "longitude";
      :units = "degrees_east";
      :valid_max = 180.0; // double
      :valid_min = -180.0; // double
      :accuracy = 0.09; // double
      :_ChunkSizes = 498U; // uint

    int longitude_qc(n_measurements=1493);
      :_FillValue = -127; // int
      :coverage_content_type = "qualityInformation";
      :long_name = "Estimated Subsurface Longitude Quality Flag";
      :standard_name = "aggregate_quality_flag";
      :valid_max = 9; // int
      :valid_min = 0; // int
      :flag_values = 1, 2, 3, 4, 9; // int
      :flag_meanings = "good not_evaluated questionable bad missing";
      :comment = "Use caution - these are estimated subsurface position values, the deviation from actual position may be several hundreds of meters! Use the gps position variables for highly accurate positions at the surface. These estimations are a dead reckoning using the GPS positions at dive start and end, and the gliders estimated velocity. The calculation methods are described in: \"Rudnick, D. L., Sherman, J. T., & Wu, A. P. (2018). Depth-average velocity from Spray underwater gliders. Journal of Atmospheric and Oceanic Technology, (2018), 35, 1665-1673; doi: https://doi.org/10.1175/JTECH-D-17-0200.1\". The accuracy attribute reflects an accuracy of approximately +/-800m (0.09 &deg; Lon)1=Good/Pass, 2=Not Evaluated, 3=Questionable, Suspect or of High Interest, 4=Fail/Bad, 9=Missing Data. See the references for more details on the flag meanings.";
      :references = "Paris. Intergovernmental Oceanographic Commission of UNESCO, 2013. Ocean Data Standards, Vol.3:Recommendation for a Quality Flag Scheme for the Exchange of Oceanographic and Marine    Meteorological Data. (IOC Manuals and Guides, 54, Vol. 3.) 12 pp. (English.)(IOC/2013/MG/54-3) https://repository.oceanbestpractices.org/bitstream/handle/11329/413/MG54_3.doc";
      :_ChunkSizes = 747U; // uint

    double pres(n_measurements=1493);
      :_FillValue = -999.0; // double
      :ancillary_variables = "pres_qc";
      :coordinates = "time longitude latitude depth";
      :coverage_content_type = "physicalMeasurement";
      :long_name = "Pressure";
      :observation_type = "measured";
      :platform = "platform_meta";
      :positive = "down";
      :reference_datum = "sea-surface";
      :sensor = "sensor_ctd";
      :standard_name = "sea_water_pressure";
      :units = "dbar";
      :valid_max = 2000.0; // double
      :valid_min = 0.0; // double
      :vocabulary = "https://vocab.nerc.ac.uk/collection/OG1/current";
      :_ChunkSizes = 498U; // uint

    int pres_qc(n_measurements=1493);
      :_FillValue = -127; // int
      :coordinates = "time longitude latitude depth";
      :coverage_content_type = "qualityInformation";
      :long_name = "Pressure Quality Flag";
      :standard_name = "aggregate_quality_flag";
      :valid_max = 9; // int
      :valid_min = 0; // int
      :flag_values = 1, 2, 3, 4, 9; // int
      :flag_meanings = "good not_evaluated questionable bad missing";
      :comment = "1=Good/Pass, 2=Not Evaluated, 3=Questionable, Suspect or of High Interest, 4=Fail/Bad, 9=Missing Data. See the references for more details on the flag meanings.";
      :references = "Paris. Intergovernmental Oceanographic Commission of UNESCO, 2013. Ocean Data Standards, Vol.3:Recommendation for a Quality Flag Scheme for the Exchange of Oceanographic and Marine    Meteorological Data. (IOC Manuals and Guides, 54, Vol. 3.) 12 pp. (English.)(IOC/2013/MG/54-3) https://repository.oceanbestpractices.org/bitstream/handle/11329/413/MG54_3.doc";
      :_ChunkSizes = 747U; // uint

    double psal(n_measurements=1493);
      :_FillValue = -999.0; // double
      :ancillary_variables = "psal_qc";
      :colorBarMaximum = 35.0; // double
      :colorBarMinimum = 32.0; // double
      :comment = "PSS-78, calculated on board glider";
      :coordinates = "time longitude latitude depth";
      :coverage_content_type = "physicalMeasurement";
      :ioos_category = "Salinity";
      :long_name = "Sea Water Practical Salinity";
      :observation_type = "measured";
      :sensor = "sensor_ctd";
      :standard_name = "sea_water_practical_salinity";
      :units = "1";
      :valid_max = 40.0; // double
      :valid_min = 0.0; // double
      :vocabulary = "https://vocab.nerc.ac.uk/collection/OG1/current";
      :_ChunkSizes = 498U; // uint

    int psal_qc(n_measurements=1493);
      :_FillValue = -127; // int
      :coverage_content_type = "qualityInformation";
      :long_name = "Sea Water Practical Salinity Quality Flag";
      :short_name = "Salinity Quality Flag";
      :valid_max = 9; // int
      :valid_min = 1; // int
      :flag_values = 1, 2, 3, 4, 9; // int
      :flag_meanings = "good not_evaluated questionable bad missing";
      :comment = "1=Good/Pass, 2=Not Evaluated, 3=Questionable, Suspect or of High Interest, 4=Fail/Bad, 9=Missing Data. See the references for more details on the flag meanings.";
      :references = "Paris. Intergovernmental Oceanographic Commission of UNESCO, 2013. Ocean Data Standards, Vol.3:Recommendation for a Quality Flag Scheme for the Exchange of Oceanographic and Marine    Meteorological Data. (IOC Manuals and Guides, 54, Vol. 3.) 12 pp. (English.)(IOC/2013/MG/54-3) https://repository.oceanbestpractices.org/bitstream/handle/11329/413/MG54_3.doc";
      :_ChunkSizes = 747U; // uint

    double temp(n_measurements=1493);
      :_FillValue = -999.0; // double
      :ancillary_variables = "temp_qc";
      :colorBarMaximum = 32.0; // double
      :colorBarMinimum = 0.0; // double
      :coordinates = "time longitude latitude depth";
      :coverage_content_type = "physicalMeasurement";
      :ioos_category = "Temperature";
      :long_name = "Sea Water Temperature";
      :sensor = "sensor_ctd";
      :observation_type = "measured";
      :standard_name = "sea_water_temperature";
      :units = "degree_C";
      :valid_max = 40.0; // double
      :valid_min = -5.0; // double
      :vocabulary = "https://vocab.nerc.ac.uk/collection/OG1/current";
      :_ChunkSizes = 498U; // uint

    int temp_qc(n_measurements=1493);
      :_FillValue = -127; // int
      :coordinates = "time longitude latitude depth";
      :coverage_content_type = "qualityInformation";
      :long_name = "Sea Water Temperature Quality Flag";
      :valid_max = 9; // int
      :valid_min = 1; // int
      :flag_values = 1, 2, 3, 4, 9; // int
      :flag_meanings = "good not_evaluated questionable bad missing";
      :comment = "1=Good/Pass, 2=Not Evaluated, 3=Questionable, Suspect or of High Interest, 4=Fail/Bad, 9=Missing Data. See the references for more details on the flag meanings.";
      :references = "Paris. Intergovernmental Oceanographic Commission of UNESCO, 2013. Ocean Data Standards, Vol.3:Recommendation for a Quality Flag Scheme for the Exchange of Oceanographic and Marine    Meteorological Data. (IOC Manuals and Guides, 54, Vol. 3.) 12 pp. (English.)(IOC/2013/MG/54-3) https://repository.oceanbestpractices.org/bitstream/handle/11329/413/MG54_3.doc";
      :_ChunkSizes = 747U; // uint

    double cndc(n_measurements=1493);
      :_FillValue = -999.0; // double
      :ancillary_variables = "psal_qc";
      :colorBarMaximum = 6.0; // double
      :colorBarMinimum = 2.0; // double
      :coordinates = "time longitude latitude depth";
      :coverage_content_type = "physicalMeasurement";
      :long_name = "Conductivity";
      :sensor = "sensor_ctd";
      :standard_name = "sea_water_electrical_conductivity";
      :ioos_category = "salinity";
      :observation_type = "calculated";
      :platform = "platform_meta";
      :units = "S m-1";
      :valid_max = 10.0; // double
      :valid_min = 0.0; // double
      :vocabulary = "https://vocab.nerc.ac.uk/collection/OG1/current";
      :_ChunkSizes = 498U; // uint

    int cndc_qc(n_measurements=1493);
      :_FillValue = -127; // int
      :comment = "1=Good/Pass, 2=Not Evaluated, 3=Questionable, Suspect or of High Interest, 4=Fail/Bad, 9=Missing Data. See the references for more details on the flag meanings.";
      :coverage_content_type = "qualityInformation";
      :long_name = "Conductivity Quality Flag";
      :valid_max = 9; // int
      :valid_min = 1; // int
      :flag_values = 1, 2, 3, 4, 9; // int
      :flag_meanings = "good not_evaluated questionable bad missing";
      :references = "Paris. Intergovernmental Oceanographic Commission of UNESCO, 2013. Ocean Data Standards, Vol.3:Recommendation for a Quality Flag Scheme for the Exchange of Oceanographic and Marine    Meteorological Data. (IOC Manuals and Guides, 54, Vol. 3.) 12 pp. (English.)(IOC/2013/MG/54-3) https://repository.oceanbestpractices.org/bitstream/handle/11329/413/MG54_3.doc";
      :_ChunkSizes = 747U; // uint

    double chla(n_measurements=1493);
      :_FillValue = -999.0; // double
      :ancillary_variables = "chla_qc";
      :comment = "Chlorophyll-a concentration estimated from fluorescence measurements. See the sensor_fchl variable for information about the fluorometer.";
      :coordinates = "time longitude latitude depth";
      :coverage_content_type = "physicalMeasurement";
      :ioos_category = "Other";
      :long_name = "Chlorophyll-a concentration";
      :observation_type = "measured";
      :sensor = "sensor_fchl";
      :standard_name = "mass_concentration_of_chlorophyll_a_in_sea_water";
      :units = "mg m-3";
      :vocabulary = "https://vocab.nerc.ac.uk/collection/OG1/current";
      :_ChunkSizes = 498U; // uint

    int chla_qc(n_measurements=1493);
      :_FillValue = -127; // int
      :coordinates = "time longitude latitude depth";
      :coverage_content_type = "qualityInformation";
      :long_name = "Chlorophyll-a concentration Quality Flag";
      :valid_max = 9; // int
      :valid_min = 1; // int
      :flag_values = 1, 2, 3, 4, 9; // int
      :flag_meanings = "good not_evaluated questionable bad missing";
      :comment = "1=Good/Pass, 2=Not Evaluated, 3=Questionable, Suspect or of High Interest, 4=Fail/Bad, 9=Missing Data. See the references for more details on the flag meanings.";
      :references = "Paris. Intergovernmental Oceanographic Commission of UNESCO, 2013. Ocean Data Standards, Vol.3:Recommendation for a Quality Flag Scheme for the Exchange of Oceanographic and Marine    Meteorological Data. (IOC Manuals and Guides, 54, Vol. 3.) 12 pp. (English.)(IOC/2013/MG/54-3) https://repository.oceanbestpractices.org/bitstream/handle/11329/413/MG54_3.doc";
      :_ChunkSizes = 747U; // uint

    double doxy(n_measurements=1493);
      :_FillValue = -999.0; // double
      :ancillary_variables = "doxy_qc";
      :coordinates = "time longitude latitude depth";
      :coverage_content_type = "physicalMeasurement";
      :ioos_category = "physical_oceanography";
      :long_name = "Dissolved Oxygen";
      :observation_type = "measured";
      :platform = "platform_meta";
      :sensor = "sensor_doxy";
      :standard_name = "moles_of_oxygen_per_unit_mass_in_sea_water";
      :units = "micromol kg-1";
      :valid_max = 500.0; // double
      :valid_min = 0.0; // double
      :vocabulary = "https://vocab.nerc.ac.uk/collection/OG1/current";
      :_ChunkSizes = 498U; // uint

    int doxy_qc(n_measurements=1493);
      :_FillValue = -127; // int
      :coordinates = "time longitude latitude depth";
      :coverage_content_type = "qualityInformation";
      :long_name = "Dissolved Oxygen Quality Flag";
      :valid_max = 9; // int
      :valid_min = 1; // int
      :flag_values = 1, 2, 3, 4, 9; // int
      :flag_meanings = "good not_evaluated questionable bad missing";
      :comment = "1=Good/Pass, 2=Not Evaluated, 3=Questionable, Suspect or of High Interest, 4=Fail/Bad, 9=Missing Data. See the references for more details on the flag meanings.";
      :references = "Paris. Intergovernmental Oceanographic Commission of UNESCO, 2013. Ocean Data Standards, Vol.3:Recommendation for a Quality Flag Scheme for the Exchange of Oceanographic and Marine    Meteorological Data. (IOC Manuals and Guides, 54, Vol. 3.) 12 pp. (English.)(IOC/2013/MG/54-3) https://repository.oceanbestpractices.org/bitstream/handle/11329/413/MG54_3.doc";
      :_ChunkSizes = 747U; // uint

    double time_gps(n_measurements=1493);
      :_FillValue = -999.0; // double
      :ancillary_variables = "gps_start_qc gps_start_qc_tests";
      :calendar = "gregorian";
      :comment = "Time from GPS at surface for the start position of the dive. These data are transmitted in near-real-time and are uncorrected. Flags are provided in the gps_start_qc and gps_start_qc_tests variables. ";
      :ioos_category = "Time";
      :long_name = "GPS Time at Dive Start";
      :observation_type = "measured";
      :platform = "platform_meta";
      :standard_name = "time";
      :units = "seconds since 1970-01-01T00:00:00Z";
      :valid_min = 1.0E9; // double
      :valid_max = 4.0E9; // double
      :_ChunkSizes = 498U; // uint

    double longitude_gps(n_measurements=1493);
      :_FillValue = -999.0; // double
      :_CoordinateAxisType = "Lon";
      :ancillary_variables = "gps_start_qc gps_start_qc_tests";
      :comment = "Longitude from GPS at surface for the starting position of the dive. These data are transmitted in near-real-time and are uncorrected. Flags are provided in the gps_end_qc and gps_end_qc_tests variables. ";
      :ioos_category = "Location";
      :long_name = "GPS Longitude at Dive Start";
      :observation_type = "measured";
      :platform = "platform_meta";
      :standard_name = "longitude";
      :units = "degrees_east";
      :valid_max = 180.0; // double
      :valid_min = -180.0; // double
      :_ChunkSizes = 498U; // uint

    double latitude_gps(n_measurements=1493);
      :_FillValue = -999.0; // double
      :ancillary_variables = "gps_start_qc gps_start_qc_tests";
      :comment = "Latitude from GPS at surface for the start position of the dive. These data are transmitted in near-real-time and are uncorrected. Flags are provided in the gps_start_qc and gps_start_qc_tests variables. ";
      :ioos_category = "Location";
      :long_name = "GPS Latitude at Dive Start";
      :observation_type = "measured";
      :platform = "platform_meta";
      :standard_name = "latitude";
      :units = "degrees_north";
      :valid_max = 90.0; // double
      :valid_min = -90.0; // double
      :_ChunkSizes = 498U; // uint

    int gps_start_qc(n_measurements=1493);
      :_FillValue = -127; // int
      :comment = "1=Good/Pass, 2=Not Evaluated, 3=Questionable, Suspect or of High Interest, 4=Fail/Bad, 9=Missing Data. See the references for more details on the flag meanings.";
      :flag_values = 1, 2, 3, 4, 9; // int
      :flag_meanings = "good not_evaluated questionable bad missing";
      :long_name = "Summary Quality Flag for the GPS Start Position";
      :references = "Paris. Intergovernmental Oceanographic Commission of UNESCO, 2013. Ocean Data Standards, Vol.3:Recommendation for a Quality Flag Scheme for the Exchange of Oceanographic and Marine    Meteorological Data. (IOC Manuals and Guides, 54, Vol. 3.) 12 pp. (English.)(IOC/2013/MG/54-3) https://repository.oceanbestpractices.org/bitstream/handle/11329/413/MG54_3.doc";
      :standard_name = "aggregate_quality_flag";
      :valid_max = 9; // int
      :valid_min = 1; // int
      :_ChunkSizes = 747U; // uint

    int gps_start_qc_tests(n_measurements=1493);
      :_FillValue = -127; // int
      :comment = "gps_good=0 gps_day_problem=1 gps_repeat=2 gps_backward=3 gps_too_fast_on_surface=4 gps_too_soon=5 gps_too_far=6 gps_bad_hdop=7 gps_bad_status=8 gps_no_surfacing=9 gps_manual=10 gps_no_dive=99";
      :long_name = "Detailed Quality Flags for the GPS Start Position";
      :flag_values = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 99; // int
      :flag_meanings = "gps_good gps_day_problem gps_repeat gps_backward gps_too_fast_on_surface gps_too_soon gps_too_far gps_bad_hdop gps_bad_status gps_no_surfacing gps_manual gps_no_dive";
      :standard_name = "quality_flag";
      :valid_max = 99; // int
      :valid_min = 0; // int
      :_ChunkSizes = 747U; // uint

    double time_gps_end(n_measurements=1493);
      :_FillValue = -999.0; // double
      :ancillary_variables = "gps_end_qc gps_end_qc_tests";
      :comment = "Time from GPS at surface for the end position of the dive. These data are transmitted in near-real-time. Flags are provided in the gps_start_qc and gps_start_qc_tests variables. This location corresponds closely with the surface value of the profile measurements.";
      :ioos_category = "Location";
      :long_name = "GPS Time at Dive End";
      :observation_type = "measured";
      :platform = "platform_meta";
      :standard_name = "time";
      :units = "seconds since 1970-01-01T00:00:00Z";
      :valid_min = 1.0E9; // double
      :valid_max = 4.0E9; // double
      :_ChunkSizes = 498U; // uint

    double latitude_gps_end(n_measurements=1493);
      :_FillValue = -999.0; // double
      :colorBarMaximum = 90.0; // double
      :colorBarMinimum = -90.0; // double
      :comment = "Latitude from GPS at surface for the end position of the dive. These data are transmitted in near-real-time. Flags are provided in the gps_start_qc and gps_start_qc_tests variables.This location corresponds closely with the surface value of the profile measurements.";
      :ioos_category = "Location";
      :long_name = "GPS Latitude at Dive End";
      :observation_type = "measured";
      :platform = "platform_meta";
      :standard_name = "latitude";
      :units = "degrees_north";
      :valid_max = 90.0; // double
      :valid_min = -90.0; // double
      :ancillary_variables = "gps_end_qc gps_end_qc_tests";
      :_ChunkSizes = 498U; // uint

    double longitude_gps_end(n_measurements=1493);
      :_FillValue = -999.0; // double
      :colorBarMaximum = 180.0; // double
      :colorBarMinimum = -180.0; // double
      :comment = "Longitude from GPS at surface for the ending position of the dive. These data are transmitted in near-real-time. Flags are provided in the gps_end_qc and gps_end_qc_tests variables. This location corresponds closely with the surface position of the profile measurements.";
      :ioos_category = "Location";
      :long_name = "GPS Longitude at Dive End";
      :observation_type = "measured";
      :platform = "platform_meta";
      :standard_name = "longitude";
      :units = "degrees_east";
      :valid_max = 180.0; // double
      :valid_min = -180.0; // double
      :ancillary_variables = "gps_end_qc gps_end_qc_tests";
      :_ChunkSizes = 498U; // uint

    int gps_end_qc(n_measurements=1493);
      :_FillValue = -127; // int
      :long_name = "Summary Quality Flag for the GPS End Postion";
      :valid_max = 9; // int
      :valid_min = 1; // int
      :flag_values = 1, 2, 3, 4, 9; // int
      :flag_meanings = "good not_evaluated questionable bad missing";
      :comment = "1=Good/Pass, 2=Not Evaluated, 3=Questionable, Suspect or of High Interest, 4=Fail/Bad, 9=Missing Data. See the references for more details on the flag meanings.";
      :references = "Paris. Intergovernmental Oceanographic Commission of UNESCO, 2013. Ocean Data Standards, Vol.3:Recommendation for a Quality Flag Scheme for the Exchange of Oceanographic and Marine    Meteorological Data. (IOC Manuals and Guides, 54, Vol. 3.) 12 pp. (English.)(IOC/2013/MG/54-3) https://repository.oceanbestpractices.org/bitstream/handle/11329/413/MG54_3.doc";
      :standard_name = "aggregate_quality_flag";
      :_ChunkSizes = 747U; // uint

    int gps_end_qc_tests(n_measurements=1493);
      :_FillValue = -127; // int
      :long_name = "Detailed Quality Flags for the GPS End Position";
      :valid_max = 99; // int
      :valid_min = 0; // int
      :flag_values = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 99; // int
      :flag_meanings = "gps_good gps_day_problem gps_repeat gps_backward gps_too_fast_on_surface gps_too_soon gps_too_far gps_bad_hdop gps_bad_status gps_no_surfacing gps_manual gps_no_dive";
      :comment = "gps_good=0 gps_day_problem=1 gps_repeat=2 gps_backward=3 gps_too_fast_on_surface=4 gps_too_soon=5 gps_too_far=6 gps_bad_hdop=7 gps_bad_status=8 gps_no_surfacing=9 gps_manual=10 gps_no_dive=99";
      :standard_name = "quality_flag";
      :_ChunkSizes = 747U; // uint

    String wmo_identifier;
      :ioos_category = "Identifier";
      :long_name = "WMO ID";

    int sensor_doxy;
      :_FillValue = -127; // int
      :_Unsigned = "false";
      :coverage_content_type = "referenceInformation";
      :ioos_category = "Identifier";
      :long_name = "Oxygen Sensor Metadata";
      :make_model = "Sea-Bird SBE 63 dissolved oxygen sensor";
      :platform = "platform_meta";
      :type = "OPTODE_DOXY";
      :type_vocabulary = "http://vocab.nerc.ac.uk/collection/R25/current/";
      :maker = "Sea-Bird Scientific";
      :maker_vocabulary = "http://vocab.nerc.ac.uk/collection/R26/current/";
      :model = "Sea-Bird SBE 63 dissolved oxygen sensor";
      :model_vocabulary = "http://vocab.nerc.ac.uk/collection/L22/current/";

    int sensor_ctd;
      :_FillValue = -127; // int
      :_Unsigned = "false";
      :coverage_content_type = "referenceInformation";
      :ioos_category = "Identifier";
      :long_name = "CTD Metadata";
      :make_model = "Sea-Bird SBE 41CP CTD";
      :platform = "platform_meta";
      :type = "CTD";
      :units = "1";
      :maker = "Sea-Bird Scientific";
      :maker_vocabulary = "https://vocab.nerc.ac.uk/collection/L35/current";
      :maker_uri = "https://vocab.nerc.ac.uk/collection/L35/current/MAN0013/";
      :model = "Sea-Bird SBE 41CP CTD";
      :model_vocabulary = "https://vocab.nerc.ac.uk/collection/L22/current";
      :model_uri = "https://vocab.nerc.ac.uk/collection/L22/current/TOOL0669/";
      :type_vocabulary = "https://vocab.nerc.ac.uk/collection/L05/current";
      :type_uri = "https://vocab.nerc.ac.uk/collection/L05/current/130/";

    int sensor_fchl;
      :_FillValue = -127; // int
      :_Unsigned = "false";
      :coverage_content_type = "referenceInformation";
      :ioos_category = "Identifier";
      :long_name = "Fluorometer Metadata";
      :platform = "platform_meta";
      :type = "fluorometer_chla";
      :type_vocabulary = "http://vocab.nerc.ac.uk/collection/R25/current/";
      :maker = "Seapoint Sensors, Inc.";
      :maker_vocabulary = "http://vocab.nerc.ac.uk/collection/R26/current/";
      :model = "Seapoint chlorophyll fluorometer";
      :model_vocabulary = "http://vocab.nerc.ac.uk/collection/L05/current";
      :model_uri = "http://vocab.nerc.ac.uk/collection/L05/current/113/";

    String platform_model;
      :ioos_category = "Identifier";
      :long_name = "Model of the glider";
      :comment = "The NERC vocabulary defines terms used to describe designs or versions of platforms.";
      :platform_model_uri = "http://vocab.nerc.ac.uk/collection/B76/current/B7600027/";
      :platform_model_vocabulary = "http://vocab.nerc.ac.uk/collection/B76/current/";

    String platform_serial_number;
      :ioos_category = "Identifier";
      :long_name = "Glider serial number";

    int platform_meta;
      :_FillValue = -127; // int
      :comment = "Spray Glider sp028";
      :coverage_content_type = "referenceInformation";
      :id = "sp028";
      :sensor = "sensor_ctd";
      :ioos_category = "Identifier";
      :long_name = "Platform Metadata";
      :platform_type = "subsurface gliders";
      :platform_type_vocabulary = "http://vocab.nerc.ac.uk/collection/L06/current/27/";
      :platform_maker = "Scripps Institution of Oceanography Instrument Development Group";
      :platform_depth_rating = "1000";
      :platform_model = "Scripps Institution of Oceanography Spray glider";
      :platform_model_uri = "http://vocab.nerc.ac.uk/collection/B76/current/B7600027/";
      :platform_model_vocabulary = "http://vocab.nerc.ac.uk/collection/B76/current/";
      :platform_serial_number = "sp028";
      :type = "platform";
      :units = "1";
      :wmo_id = "4801921";
      :wmo_identifier = "4801921";

    double deployment_time(n_measurements=1493);
      :_FillValue = -999.0; // double
      :comment = "GPS Time value for the start position of the first dive.";
      :ioos_category = "Location";
      :long_name = "Deployment Time, GPS at start of first dive";
      :observation_type = "measured";
      :platform = "platform_meta";
      :standard_name = "time";
      :units = "seconds since 1970-01-01T00:00:00Z";
      :_ChunkSizes = 498U; // uint

    double deployment_latitude(n_measurements=1493);
      :_FillValue = -999.0; // double
      :comment = "GPS latitude value for the start position of the first dive.";
      :ioos_category = "Location";
      :long_name = "Deployment Latitude, GPS at start of first dive";
      :observation_type = "measured";
      :platform = "platform_meta";
      :standard_name = "latitude";
      :units = "degrees_north";
      :_ChunkSizes = 498U; // uint

    double deployment_longitude(n_measurements=1493);
      :_FillValue = -999.0; // double
      :comment = "GPS longitude value for the start position of the first dive.";
      :ioos_category = "Location";
      :long_name = "Deployment longitude, GPS at start of first dive";
      :observation_type = "measured";
      :platform = "platform_meta";
      :standard_name = "longitude";
      :units = "degrees_east";
      :_ChunkSizes = 498U; // uint

  // global attributes:
  :Conventions = "CF-1.10, ACDD-1.3, OG-1.0";
  :acknowledgement = "Funded by National Oceanic and Atmospheric Administration (NOAA): Global Ocean Monitoring and Observing (GOMO) Program and Integrated Ocean Observing System. Supported by Instrument Development Group - Scripps Institution of Oceanography";
  :cdm_trajectory_variables = "trajectory";
  :comment = "This file contains data from the following specific sensors: Sea-Bird SBE 41CP CTD, Seapoint chlorophyll fluorometer, Sea-Bird SBE 63 dissolved oxygen sensor.";
  :contributing_institutions = "Scripps Institution of Oceanography";
  :contributing_institutions_role = "Operator";
  :contributing_institutions_vocabulary = "https://vocab.nerc.ac.uk/collection/W08/current/";
  :contributor_email = "drudnick@ucsd.edu, jpsevadjian@ucsd.edu";
  :contributor_name = "Daniel Rudnick, Jennifer Sevadjian";
  :contributor_role = "principalInvestigator, resourceProvider";
  :contributor_role_vocabulary = "https://vocab.nerc.ac.uk/collection/G04/current";
  :creator_email = "idgdata@ucsd.edu";
  :creator_institution = "Scripps Institution of Oceanography";
  :creator_name = "Instrument Development Group";
  :creator_type = "group";
  :creator_url = "https://spraydata.ucsd.edu";
  :data_url = "https://spraydata.ucsd.edu/erddap/info/sp028_20230202T1637_R/index.html";
  :date_created = "2024-05-31T20:07:33Z";
  :date_issued = "2024-05-31T20:07:33Z";
  :date_metadata_modified = "2024-05-31T20:07:33Z";
  :date_modified = "2024-05-31T20:07:33Z";
  :doi = "10.21238/S8SPRAY1618";
  :featureType = "trajectory";
  :geospatial_bounds = "POLYGON ((-123.5721 38.318775, -123.0713 38.318775, -123.0713 38.2429, -123.5721 38.2429, -123.5721 38.318775))";
  :geospatial_bounds_crs = "EPSG:4326";
  :geospatial_lat_max = 38.318775; // double
  :geospatial_lat_min = 38.2429; // double
  :geospatial_lat_units = "degrees_north";
  :geospatial_lon_max = -123.0713; // double
  :geospatial_lon_min = -123.5721; // double
  :geospatial_lon_units = "degrees_east";
  :geospatial_vertical_max = 0.03969955209296338; // double
  :geospatial_vertical_min = 501.6665808273762; // double
  :geospatial_vertical_positive = "down";
  :geospatial_vertical_units = "EPSG:5831";
  :history = "2023-06-16T15:40:09Z: Jenn readsat(maxdives=3000, Gps_Good=0, Gps_Bad=8, Gps_No_Dive=99, Gps_No_Surfacing=9, DOConv=44660). \n2023-06-16T15:40:49Z: Jenn fixgps3(R=6378000, Too_Soon=60, Too_Fast_On_Surface=5, Too_Far=100, Bad_HDOP=12, Gps_Good=0, Gps_Repeat=2, Gps_Backward=3, Gps_Too_Fast_On_Surface=4, Gps_Too_Soon=5, Gps_Too_Far=6, Gps_Bad_HDOP=7, Gps_Bad_Status=8, Gps_No_Surfacing=9). \n2023-06-16T15:40:49Z: Jenn calcvelsat(R=6378000, Gps_No_Surfacing=9). \n2023-06-16T15:42:15Z: Jenn calox(filename=/Users/Shared/spray/data/ox/doxcal.xlsx, sheetname=AllOxMissions, DOConv=44660, Gain=1.0811, Offset=-0.0615). \n;2024-05-31T20:07:33Z: OG-1.0 NetCDF created by J.P. Sevadjian with make_mission_nc_og10.py, input file: 23202801_aug.mat, with MD5 checksum: b0936e175fd11895c04fdba38f379df0, output file: ./mission_output/OG-10-202400415/sp028_20230202T1637_R.nc.";
  :id = "sp028-20230202T1637";
  :infoUrl = "https://spraydata.ucsd.edu";
  :institution = "Scripps Institution of Oceanography";
  :instrument = "This file contains data from the following specific sensors: Sea-Bird SBE 41CP CTD, Seapoint chlorophyll fluorometer, Sea-Bird SBE 63 dissolved oxygen sensor.";
  :internal_mission_identifier = "23202801";
  :keywords = "AUVS > Autonomous Underwater Vehicles, Earth Science > Oceans > Ocean Pressure > Water Pressure, Earth Science > Oceans > Ocean Temperature > Water Temperature, Earth Science > Oceans > Salinity/Density > Conductivity, Earth Science > Oceans > Salinity/Density > Density, Earth Science > Oceans > Salinity/Density > Salinity, glider, In Situ Ocean-based platforms > Seaglider, Slocum, Spray, trajectory, underwater glider, water, wmo, underwater glider, pressure, temperature, salinity, currents, oxygen, fluorescence, chlorophyll;";
  :keywords_vocabulary = "GCMD Science Keywords";
  :license = "The data may be used and redistributed for free but is not intended for legal use, since it may contain inaccuracies. Neither the data Contributor, University of California, IOOS, NOAA, nor the United States Government, nor any of their employees or contractors, makes any warranty, express or implied, including warranties of merchantability and fitness for a particular purpose, or assumes any legal liability for the accuracy, completeness, or usefulness, of this information.";
  :metadata_link = "https://spraydata.ucsd.edu";
  :mission_id = "23202801";
  :naming_authority = "edu.ucsd.idg";
  :network = "OceanGliders > BOON > Northeast Pacific Ocean > California Underwater Glider Network, California Underwater Glider Network (CUGN), IOOS";
  :platform = "sub-surface gliders";
  :platform_institution = "Scripps Institution of Oceanography";
  :platform_type = "Spray Glider";
  :platform_vocabulary = "https://vocab.nerc.ac.uk/collection/L06/current/";
  :processing_level = "This is a near-real-time data product. Within the Spray program to is considered a Level 2 product. Real-time quality control has been conducted and users should apply the supplied QARTOD flags. Afer a mission is complete a higher-quality data product is provided at https://spraydata.ucsd.edu and should be used in place of the near-real-time data as soon as it is available.";
  :project = "California Underwater Glider Network (CUGN)";
  :publisher_email = "idgdata@ucsd.edu";
  :publisher_institution = "University of California - San Diego; Scripps Institution of Oceanography";
  :publisher_name = "Instrument Development Group";
  :publisher_type = "group";
  :publisher_url = "https://spraydata.ucsd.edu";
  :references = "Rudnick, D. L. (2016). Ocean research enabled by underwater gliders. Annual review of marine science, 8, 519-541, doi:10.1146/annurev-marine-122414-033913\n Rudnick, D. L., Davis, R. E., & Sherman, J. T. (2016). Spray Underwater Glider Operations. Journal of Atmospheric and Oceanic Technology, 33(6), 1113-1122, doi:10.1175/JTECH-D-15-0252.1\n Rudnick, D. L., Davis, R. E., Eriksen, C. C., Fratantoni, D. M., & Perry, M. J. (2004). Underwater gliders for ocean research. Marine Technology Society Journal, 38(2), 73-84, doi:10.4031/002533204787522703\n Sherman, J., Davis, R. E., Owens, W. B., & Valdes, J. (2001). The autonomous underwater glider \'Spray\'. IEEE Journal of oceanic Engineering, 26(4), 437-446, doi:10.1109/48.972076";
  :rtqc_method = "Spray Data Center RTQC";
  :sea_name = "Coastal Waters of California";
  :site = "CUGN Line 56";
  :source = "Spray Underwater Glider";
  :standard_name_vocabulary = "CF Standard Name Table v83";
  :summary = "Spray glider data from mission 23202801, part of the California Underwater Glider Network (CUGN) project. This is the near-real-time dataset for the full mission, spanning from 2023-02-02 to 2023-05-25. \n\nThe overarching goal of the California Underwater Glider Network is to sustain baseline observations of climate variability off the coast of California. The technical approach is to deploy autonomous underwater gliders in a network to provide real-time data.\nThe CUGN uses Spray underwater gliders making repeated dives from the surface to 500 m and back, repeating the cycle every 3 hours, and traveling 3 km in the horizontal during that time. The CUGN includes gliders on three of the traditional cross-shore CalCOFI lines: line 66.7 off Monterey Bay, line 80 off Point Conception, and line 90 off Dana Point.\n The glider missions typically last about 100 days, and cover over 2000 km, thus providing 4-6 sections on lines extending 300-500 km offshore. Since 2005 the CUGN has covered 200,000 km over ground in 28 glider-years, while doing 90,000 dives.";
  :time_coverage_duration = "P0000-03-22T21:25:00";
  :time_coverage_end = "2023-05-25T14:02:00Z";
  :time_coverage_resolution = "P0000-00-00T00:00:04";
  :time_coverage_start = "2023-02-02T16:37:00Z";
  :title = "Near-real-time Data from Spray Glider Mission 23202801 (sp028-20230202T1637)";

  data:
    trajectory =   "sp028-20230202T1637"
    profile_index = 
      {2, 3, 4, 5, 6, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50}
    time_profile = 
      {1.675361294999998E9, 1.6753642950000005E9, 1.6753672950000026E9, 1.6753702949999971E9, 1.675373415E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9}
    time_profile_qc = 
      {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
    latitude_profile = 
      {38.3187, 38.3187, 38.318775, 38.3187, 38.3187, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735}
    latitude_profile_qc = 
      {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
    latitude_uv = 
      {38.3187, 38.3187, 38.31875, 38.3187, 38.3187, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.253, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2513, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2436, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2426, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.2442, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24535, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24555, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24625, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.24685, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.2474, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.24875, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.25, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2495, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.2483, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.24635, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.2551, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28, 38.28}
    latitude_uv_qc = 
      {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
    longitude_profile = 
      {-123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721}
    longitude_profile_qc = 
      {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
    longitude_uv = 
      {-123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.3425, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35065, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.35855, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.366, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.373, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.37985, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3876, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.3961, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.40485, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4136, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.4229, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.433, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.44675, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.4647, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.48405, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.50575, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5308, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.5521, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568, -123.568}
    longitude_uv_qc = 
      {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
    time_uv = 
      {1.6753605899999974E9, 1.6753635899999995E9, 1.675366590000002E9, 1.675369589999999E9, 1.6753727099999993E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.675447590000002E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754504400000029E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754531700000012E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754558999999995E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754586299999976E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.6754616000000017E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.675464990000001E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.67546838E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.6754719500000033E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675475940000002E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.675480139999998E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754843699999971E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.6754892600000026E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.67549487E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.675500959999999E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755076199999995E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755147600000014E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755222900000002E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9, 1.6755305699999995E9}
    time_uv_qc = 
      {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
    time = 
      {1.675361294999998E9, 1.6753642950000005E9, 1.6753672950000026E9, 1.6753702949999971E9, 1.675373415E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.6754482950000026E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.675451070000003E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754538150000005E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754565299999995E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754592449999986E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754623800000029E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754658149999995E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754691600000012E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754728650000043E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754769300000007E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754811299999993E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.6754853749999976E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675490580000002E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.675496265E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755024599999979E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755093E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.6755165600000024E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.675524135000001E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9, 1.6755327749999988E9}
    time_qc = 
      {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
    wcur_x = 
      {0.0011, 7.0E-4, 0.0011, 0.0014, 0.0011, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0735, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0528, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0468, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0242, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0088, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0057, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0024, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, -0.0051, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0332, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0477, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0395, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.0305, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0029, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0086, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0097, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0216, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0604, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703, -0.0703}
    wcur_y = 
      {7.0E-4, 4.0E-4, 0.0043, 7.0E-4, 7.0E-4, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1443, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1299, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1411, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1603, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.1739, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0976, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0774, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.0922, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.1006, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0878, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0926, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0695, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0308, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0073, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, -0.0036, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0078, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0135, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.0398, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069, 0.069}
    wcur_qc = 
      {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
    wcur_qc_tests = 
      {0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0}
    depth = 
      {0.0397, 0.0794, 0.0794, 0.0397, 0.0397, 111.3673, 111.0896, 110.3754, 109.9786, 109.066, 108.4708, 107.5979, 106.8836, 105.8916, 105.3361, 104.0664, 103.2728, 102.2411, 101.4078, 100.1778, 99.3445, 97.4398, 96.0906, 94.305, 92.8764, 91.6066, 90.2177, 88.9479, 87.6384, 85.8923, 84.5828, 83.3923, 81.9637, 80.6144, 79.5032, 78.1143, 76.9634, 75.8919, 74.5426, 73.3918, 72.3599, 70.9312, 69.701, 68.7088, 67.5579, 65.9704, 64.8195, 63.7876, 62.5176, 61.4461, 60.4935, 59.3029, 58.271, 57.3582, 56.4056, 55.1356, 54.064, 53.1511, 51.9604, 50.5713, 49.4203, 48.428, 47.0785, 46.0069, 45.0146, 43.943, 42.4744, 41.2042, 40.1326, 38.267, 36.9969, 35.8458, 34.2977, 32.9482, 31.8764, 30.3284, 29.1376, 27.9864, 26.5574, 25.4063, 24.3345, 23.0246, 21.9528, 21.0001, 19.6108, 18.4596, 17.229, 16.1572, 14.8075, 13.696, 12.8226, 11.7111, 10.7187, 9.2101, 8.1383, 6.9473, 5.9946, 5.0815, 3.8111, 2.9378, 1.9056, 108.5105, 108.1137, 107.3201, 106.5662, 105.7726, 105.0584, 104.3442, 103.3522, 102.5586, 101.6856, 100.7333, 99.781, 98.9477, 97.8366, 96.924, 95.8922, 94.9399, 93.2336, 92.0431, 90.4558, 89.2257, 88.0352, 86.8447, 85.6542, 84.305, 83.1145, 81.4478, 80.0588, 78.8286, 77.1222, 75.7729, 73.9474, 72.6774, 71.3281, 69.7407, 68.3119, 67.161, 65.4942, 64.1448, 62.9939, 61.5254, 60.2951, 59.2632, 57.8741, 56.8025, 55.8103, 54.5799, 53.5083, 52.6352, 51.3254, 50.2141, 49.1821, 48.0311, 46.6816, 45.4115, 44.2605, 42.6728, 41.3233, 40.2119, 38.6639, 37.3144, 36.0442, 34.4168, 33.0276, 31.9161, 30.2093, 28.9391, 27.9071, 26.4384, 25.2475, 24.2551, 22.8658, 21.7146, 20.6825, 19.3329, 18.142, 17.0702, 15.8396, 14.3708, 13.2196, 12.1081, 10.4805, 9.3689, 7.9398, 6.5901, 5.3991, 4.4066, 3.0172, 1.8659, 110.6531, 110.3754, 109.8199, 109.2644, 108.7089, 107.9947, 107.3995, 106.6059, 105.8917, 105.1775, 104.2648, 103.3919, 102.5586, 101.5269, 100.5746, 99.5826, 98.6302, 96.6065, 95.297, 93.5511, 92.1225, 90.9717, 89.5035, 88.3924, 87.0035, 85.1781, 83.9082, 82.678, 81.17, 79.8207, 78.6699, 77.2016, 75.892, 74.7411, 73.1537, 71.725, 70.4947, 68.6295, 67.2007, 65.2561, 63.7083, 62.4383, 60.6523, 59.2632, 57.6757, 56.3263, 55.1753, 53.7465, 52.4367, 51.2857, 49.8569, 48.6265, 47.4755, 45.9275, 44.578, 43.3873, 41.7996, 40.4898, 39.4181, 37.9495, 36.8381, 35.687, 34.1787, 33.0276, 31.8765, 30.3681, 29.1773, 27.9071, 26.5971, 25.0887, 23.8979, 22.3895, 21.1589, 20.0871, 18.7771, 17.626, 16.6335, 15.4029, 14.0532, 12.8226, 11.7508, 10.0835, 8.5353, 7.3443, 6.1137, 4.9624, 3.9699, 2.6599, 1.5086, 108.4312, 108.0741, 107.4392, 106.844, 106.0504, 105.4156, 104.5823, 103.9077, 103.1538, 102.3205, 101.4476, 100.6143, 99.7413, 98.8287, 97.797, 96.924, 95.8129, 94.2257, 93.1543, 91.7257, 90.6543, 89.6622, 88.5511, 87.5591, 86.4083, 85.2971, 84.0273, 82.6383, 81.4081, 80.2176, 78.7493, 77.4397, 76.2888, 74.3442, 72.9553, 71.2488, 69.8994, 68.6692, 67.042, 65.653, 64.4623, 62.6764, 61.327, 60.057, 58.5092, 57.1201, 55.8897, 54.3021, 52.8733, 51.3651, 50.0553, 48.8646, 47.3564, 46.1657, 45.1337, 43.4667, 42.3553, 41.2836, 39.9341, 38.8227, 37.8304, 36.719, 35.4489, 34.3772, 33.4642, 32.0352, 30.8841, 29.8521, 28.8597, 27.4704, 26.359, 25.3666, 24.0964, 22.9849, 22.0322, 20.9207, 19.7299, 18.6581, 17.7054, 16.4351, 15.3236, 14.212, 13.2196, 11.9096, 10.7981, 9.885, 7.4237, 6.4313, 5.3594, 4.089, 3.0569, 2.0644, 1.0322, 106.6853, 106.3679, 105.8124, 104.9394, 104.1855, 103.511, 102.5983, 101.7254, 100.9715, 99.9794, 99.0271, 98.0748, 97.1621, 96.051, 95.2971, 94.2257, 93.0749, 91.5273, 90.2972, 88.6702, 87.44, 86.4083, 85.2178, 84.1463, 82.9558, 81.7653, 80.3764, 79.1461, 78.035, 76.5666, 75.257, 74.2252, 72.7172, 71.5663, 70.336, 68.9867, 67.7961, 66.7245, 65.4545, 64.0655, 62.7558, 61.5652, 60.057, 58.787, 57.6757, 56.0882, 54.7387, 53.5084, 51.8414, 50.4919, 49.3012, 47.6342, 46.3245, 44.8162, 43.5064, 42.395, 40.9661, 39.7754, 38.7037, 37.3144, 36.0443, 35.0123, 33.8215, 32.5116, 31.3208, 30.249, 28.7407, 27.5498, 26.5972, 25.2475, 24.1758, 23.3025, 22.1513, 20.762, 19.7299, 18.8169, 17.626, 16.5939, 15.6808, 14.609, 13.2593, 12.2272, 11.1156, 10.0438, 7.6619, 6.5504, 5.3594, 4.3272, 3.3348, 2.2629, 1.1116, 154.8105, 153.7791, 152.47, 151.0418, 149.574, 147.9475, 146.0433, 144.0993, 141.7984, 138.6246, 135.6887, 133.0306, 130.0153, 126.762, 123.6673, 120.5329, 117.3191, 113.8274, 110.6135, 107.717, 104.6617, 101.8047, 98.67, 95.813, 92.8765, 90.0988, 86.9242, 84.0273, 81.051, 78.2334, 75.2967, 72.5981, 69.8598, 67.3198, 64.8195, 62.2002, 59.6601, 57.0407, 54.2228, 51.2857, 48.6265, 45.9275, 43.5064, 41.1249, 38.5449, 36.2427, 33.6627, 31.3605, 28.9391, 26.3193, 23.8185, 21.3177, 18.8169, 16.5939, 13.9342, 11.6317, 9.0911, 6.3519, 4.1287, 1.8659, 162.5063, 161.3162, 160.0468, 158.5791, 157.1906, 155.5245, 153.66, 151.7955, 149.4153, 146.0829, 142.8298, 139.9337, 136.5615, 133.1496, 129.8169, 126.9207, 123.945, 120.9296, 118.1126, 115.2161, 112.161, 109.4628, 106.606, 103.9078, 101.0111, 98.3525, 95.6542, 92.9162, 90.3765, 87.7575, 85.0987, 82.5987, 79.9001, 77.0032, 74.2252, 71.2488, 68.1929, 65.0973, 62.3192, 59.5808, 56.7232, 54.064, 51.127, 48.5471, 45.9275, 43.5461, 41.2043, 38.8624, 36.719, 34.4565, 32.4322, 29.9315, 27.5498, 25.0887, 22.6673, 20.2459, 17.7847, 15.5617, 13.2196, 10.9966, 8.4559, 6.1137, 3.9699, 1.8659, 149.2566, 148.0268, 146.5986, 145.0514, 143.4249, 141.719, 140.0131, 138.0294, 135.5697, 132.4751, 129.7376, 127.2777, 124.7782, 121.9612, 119.1442, 116.5652, 113.9861, 111.2484, 108.7089, 106.1298, 103.3919, 100.9317, 98.3128, 95.6145, 92.6384, 89.9797, 87.2019, 84.7812, 82.2415, 79.662, 77.4, 74.8205, 72.36, 69.8201, 67.1214, 64.5417, 61.843, 59.0648, 56.485, 53.8259, 51.127, 48.6265, 46.2848, 43.8239, 41.4821, 38.9021, 36.4809, 34.1787, 31.8368, 29.4948, 27.272, 24.9697, 22.5483, 20.0474, 17.745, 15.4029, 12.9814, 10.679, 7.2252, 5.0418, 2.779, 0.9925, 181.6255, 180.4356, 179.0473, 177.54, 175.9137, 174.2874, 172.4628, 170.5588, 168.2581, 165.283, 162.5459, 160.1261, 157.746, 155.0088, 152.5889, 150.0897, 147.5507, 145.0911, 142.5521, 139.9337, 137.3947, 134.7762, 132.1577, 129.6979, 127.1984, 124.6195, 122.1596, 119.4219, 116.9619, 114.4226, 111.7245, 109.2247, 106.6456, 104.0268, 101.5666, 99.1461, 96.5272, 94.1066, 91.7654, 89.4241, 87.1226, 84.5828, 82.2415, 79.7811, 77.2809, 74.7411, 72.1219, 69.6613, 67.042, 64.3433, 61.8033, 59.2236, 56.6438, 54.3418, 52.0002, 49.5791, 47.1579, 44.578, 42.1966, 39.815, 37.4335, 35.4092, 33.1864, 31.2414, 28.82, 26.5971, 24.3345, 22.0719, 19.7696, 17.3878, 15.3236, 12.8226, 10.5996, 8.0192, 5.7961, 3.8111, 1.985, 205.9781, 204.9073, 203.5589, 202.1311, 200.5843, 198.9582, 197.2131, 195.3887, 193.2866, 190.5498, 187.8924, 185.5126, 183.0534, 180.2769, 177.6193, 174.8427, 171.9471, 168.8927, 166.1557, 163.2996, 160.3245, 157.627, 154.8898, 152.1525, 149.3359, 146.678, 143.9803, 141.2032, 138.5055, 135.6887, 132.8322, 130.2137, 127.5555, 124.8575, 122.3183, 119.779, 117.2, 114.7797, 112.2403, 109.5818, 106.963, 104.2252, 101.4476, 98.8287, 96.2494, 93.5114, 91.0511, 88.6305, 86.0908, 83.9082, 81.4081, 79.1064, 76.6857, 74.1061, 71.725, 68.7882, 65.8514, 63.2717, 60.6126, 57.9535, 55.5325, 53.0321, 50.4126, 48.1899, 45.8481, 43.5858, 41.1249, 38.4655, 36.2427, 33.5833, 31.0429, 28.6216, 26.2796, 23.9773, 21.6749, 19.2535, 16.9511, 14.5296, 12.3066, 9.885, 7.5031, 5.3594, 3.0172, 1.5483, 207.4852, 206.2557, 204.7883, 203.2019, 201.6155, 199.9101, 198.0856, 196.0629, 193.6832, 190.9068, 188.3684, 186.1869, 183.9657, 181.4272, 178.9679, 176.469, 173.9304, 171.2727, 168.5357, 165.997, 163.4186, 160.6815, 158.103, 155.4451, 152.6682, 150.1293, 147.4714, 144.6547, 142.0363, 139.1006, 136.3235, 133.5066, 130.7691, 127.9125, 124.8972, 122.1596, 119.2235, 116.4461, 113.7084, 111.169, 108.4708, 105.6933, 103.0745, 100.3762, 97.7176, 95.2971, 92.8368, 90.2178, 87.7575, 85.0987, 82.4399, 80.0192, 77.2016, 74.4236, 71.5662, 68.8676, 65.9705, 63.232, 60.5333, 57.7551, 55.215, 52.7146, 50.0553, 47.6739, 45.2131, 42.6332, 40.1723, 37.5923, 35.0122, 32.4322, 29.8521, 27.5895, 25.446, 23.1834, 21.1192, 18.7375, 16.5938, 14.4105, 12.2669, 9.8453, 7.384, 5.1609, 2.8187, 1.3101, 206.1368, 204.9073, 203.4795, 201.9328, 200.3463, 198.5616, 196.7768, 194.754, 192.3346, 189.5979, 187.1784, 184.9573, 182.7757, 180.2372, 177.9763, 175.279, 172.7404, 170.1224, 167.544, 165.045, 162.3872, 159.9278, 157.3493, 154.6517, 151.9542, 149.4946, 146.9953, 144.3373, 141.6793, 139.0609, 136.3631, 133.943, 131.3245, 128.6663, 126.3652, 123.7863, 121.4057, 118.8664, 116.2874, 113.9068, 111.6054, 109.3834, 106.9234, 104.4236, 101.8444, 99.1461, 96.4478, 93.9479, 91.4082, 88.7495, 86.3289, 83.9082, 81.4875, 79.1064, 76.6857, 74.4236, 72.1615, 69.7804, 67.3992, 64.8592, 62.3986, 59.7792, 57.1201, 54.6593, 52.1589, 49.6584, 47.277, 44.8559, 42.6332, 40.331, 38.1083, 35.7664, 33.3451, 31.0826, 28.7803, 26.5178, 24.1758, 21.6353, 19.452, 16.9908, 14.8075, 12.5051, 10.1232, 7.5825, 5.28, 3.2157, 1.5086, 293.6475, 291.2689, 288.3353, 284.7673, 279.6927, 273.6664, 267.8779, 262.0892, 256.5383, 250.9079, 245.2773, 239.5673, 233.8571, 228.0675, 222.1984, 216.567, 210.6976, 205.2245, 199.7514, 194.4367, 188.8839, 183.2517, 177.4606, 171.7487, 166.1953, 160.8798, 155.7228, 150.8037, 145.7258, 140.6478, 135.4903, 130.412, 125.1749, 119.779, 113.9861, 108.1137, 102.5586, 97.1621, 92.3209, 87.4003, 82.4796, 77.0825, 72.0028, 67.161, 62.1605, 57.3979, 52.8733, 47.9517, 43.0301, 37.9495, 33.0276, 28.3437, 23.8185, 19.2932, 14.6884, 9.7659, 5.1609, 1.985, 309.7419, 306.8878, 303.558, 299.7524, 294.8368, 289.0488, 283.4193, 277.4725, 271.4462, 264.9439, 258.2829, 251.8595, 245.9117, 239.9638, 234.2536, 228.5433, 222.8328, 217.3602, 211.8873, 206.4143, 200.9015, 195.2696, 189.8755, 184.4813, 179.2455, 173.9303, 168.2977, 162.2682, 156.7145, 151.2401, 146.0035, 140.9255, 135.9267, 131.0071, 126.1668, 121.3263, 116.3271, 111.169, 106.0901, 100.9317, 96.051, 91.0511, 85.813, 80.416, 75.3364, 70.336, 64.9386, 59.7792, 55.1753, 50.2538, 45.2528, 40.1723, 34.7741, 29.5345, 24.4536, 19.6902, 14.8472, 10.2423, 5.3991, 2.1438, 332.0976, 329.2438, 326.1522, 322.5056, 317.749, 312.5167, 307.6806, 302.6859, 297.4532, 292.2203, 286.9081, 281.3578, 275.9659, 270.6532, 265.1025, 259.631, 254.1592, 248.6874, 243.374, 237.9812, 232.7864, 227.4726, 222.0794, 217.0032, 212.0063, 207.0092, 202.0914, 197.1734, 192.176, 187.0991, 181.9428, 176.707, 171.471, 166.1557, 160.9988, 155.9212, 150.9227, 145.8448, 141.0842, 136.1647, 131.1658, 126.0874, 121.1676, 116.1684, 111.169, 106.4075, 101.9634, 97.5192, 92.9161, 88.3924, 83.7891, 79.027, 73.9474, 69.1851, 64.2639, 59.5807, 55.0562, 50.611, 46.1657, 41.3233, 36.4015, 31.5192, 26.9544, 22.6276, 18.2214, 13.7754, 9.0911, 4.5654, 1.9056, 371.135, 368.8366, 365.9041, 362.3374, 357.5818, 352.509, 347.9117, 343.0764, 338.0033, 333.1678, 328.6493, 323.9722, 319.295, 314.6969, 309.8609, 304.7076, 299.6335, 294.48, 289.2471, 283.9347, 278.5033, 272.9528, 267.7193, 262.4857, 257.3313, 252.256, 247.4186, 242.4224, 237.5846, 232.7468, 228.0675, 223.5467, 219.1051, 214.6634, 210.2217, 205.3832, 200.6239, 195.7059, 190.8671, 186.0282, 181.1098, 176.2707, 171.4314, 166.4333, 161.5938, 156.6749, 151.9145, 146.9953, 142.1554, 137.1566, 131.999, 126.9206, 122.0008, 117.0809, 112.0816, 107.0027, 102.0824, 97.4795, 93.0352, 88.3527, 83.6304, 79.1858, 74.5427, 70.0185, 65.4942, 60.9301, 56.5247, 52.278, 47.793, 43.1888, 38.6243, 34.3375, 30.1299, 25.962, 21.7146, 17.3878, 12.9814, 8.5353, 4.486, 1.8659, 403.6672, 401.1314, 398.1994, 394.871, 390.2746, 385.5196, 381.0815, 376.0886, 370.8577, 365.706, 360.6334, 355.7192, 350.8842, 346.1283, 341.293, 336.2991, 330.9879, 325.8352, 320.7616, 315.6086, 310.733, 305.8176, 300.9021, 295.9865, 290.8329, 285.8378, 280.8425, 275.9264, 270.8516, 265.7766, 260.9395, 256.0229, 251.1855, 246.5066, 241.9069, 237.3864, 232.8658, 228.2658, 223.5071, 218.9069, 214.1876, 209.5079, 204.6694, 199.8308, 195.1507, 190.5499, 185.7902, 181.0305, 176.35, 171.5901, 166.9094, 162.3079, 157.5476, 152.946, 148.3442, 143.7423, 139.0609, 134.3795, 129.5392, 124.4608, 119.3822, 114.3036, 109.066, 104.0665, 99.3048, 94.4638, 89.5432, 84.5431, 79.543, 74.7808, 69.7804, 64.7798, 60.2554, 55.731, 51.4445, 46.761, 41.9981, 37.3144, 32.6306, 28.2643, 23.9376, 19.6505, 15.2045, 10.7584, 6.3519, 2.6996, 402.4781, 399.6252, 396.2969, 392.4931, 387.5796, 382.4283, 377.7524, 372.9971, 368.1625, 363.4863, 358.8892, 354.292, 349.774, 345.0974, 340.4999, 335.7437, 331.146, 326.3897, 321.7125, 317.1145, 312.3975, 307.5614, 302.8045, 297.9682, 293.2111, 288.2953, 283.4587, 278.3841, 273.3093, 268.1552, 263.0009, 257.9258, 252.6919, 247.6958, 242.6997, 237.7033, 232.6276, 227.5517, 222.3964, 217.3203, 212.2837, 207.2073, 202.0515, 196.9749, 191.9775, 187.1386, 182.3789, 177.5398, 172.8592, 168.2579, 163.7358, 159.1342, 154.5326, 149.8515, 145.2496, 140.8063, 136.0456, 131.6021, 127.4759, 123.0323, 118.0727, 113.2321, 108.3517, 103.4711, 98.5508, 93.8287, 89.4637, 85.0192, 80.654, 76.2887, 71.8043, 67.5578, 63.232, 58.9457, 54.7783, 50.4919, 46.3641, 42.1568, 37.6319, 33.1069, 28.82, 24.3742, 20.1665, 15.9587, 11.9096, 6.5901, 2.5408, 501.6666, 497.627, 492.6369, 485.5872, 478.5372, 470.9324, 463.169, 455.4844, 447.7996, 440.1937, 432.5876, 424.9019, 416.7405, 408.8165, 401.0507, 393.2053, 385.2804, 377.4345, 369.5882, 361.9002, 354.0534, 346.2062, 338.5966, 331.1452, 323.9314, 316.7966, 309.5823, 302.5263, 295.3908, 288.0964, 280.8018, 273.5862, 266.4497, 259.2336, 252.0965, 244.642, 237.4252, 230.1288, 222.9114, 215.9317, 209.0708, 202.17, 195.1896, 188.209, 181.0695, 174.0884, 167.0278, 160.2049, 153.4611, 146.5584, 139.5761, 132.911, 125.9283, 118.7866, 111.5654, 104.1851, 96.9633, 89.8206, 82.6777, 75.6139, 68.4308, 61.5252, 54.937, 48.5072, 42.1567, 36.0441, 29.7726, 23.5009, 17.9435, 12.2271, 6.5106, 2.0644}
    depth_qc = 
      {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
    latitude = 
      {38.3187, 38.3187, 38.318775, 38.3187, 38.3187, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25265, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.25105, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.2491, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.246275, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.2429, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.24305, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.2447, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245425, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246525, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.246925, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.2477, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.249225, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.2501, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24925, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.24805, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.245675, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.2603, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735, 38.28735}
    latitude_qc = 
      {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
    longitude = 
      {-123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.3446, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.352475, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.360425, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.36765, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.3746, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.381525, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.38955, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.39815, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.407025, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.4159, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.42545, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.4356, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.451125, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.46945, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.489425, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.511725, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.53755, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5559, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721, -123.5721}
    longitude_qc = 
      {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
    pres = 
      {0.04, 0.08, 0.08, 0.04, 0.04, 112.24, 111.96, 111.24, 110.84, 109.92, 109.32, 108.44, 107.72, 106.72, 106.16, 104.88, 104.08, 103.04, 102.2, 100.96, 100.12, 98.2, 96.84, 95.04, 93.6, 92.32, 90.92, 89.64, 88.32, 86.56, 85.24, 84.04, 82.6, 81.24, 80.12, 78.72, 77.56, 76.48, 75.12, 73.96, 72.92, 71.48, 70.24, 69.24, 68.08, 66.48, 65.32, 64.28, 63.0, 61.92, 60.96, 59.76, 58.72, 57.8, 56.84, 55.56, 54.48, 53.56, 52.36, 50.96, 49.8, 48.8, 47.44, 46.36, 45.36, 44.28, 42.8, 41.52, 40.44, 38.56, 37.28, 36.12, 34.56, 33.2, 32.12, 30.56, 29.36, 28.2, 26.76, 25.6, 24.52, 23.2, 22.12, 21.16, 19.76, 18.6, 17.36, 16.28, 14.92, 13.8, 12.92, 11.8, 10.8, 9.28, 8.2, 7.0, 6.04, 5.12, 3.84, 2.96, 1.92, 109.36, 108.96, 108.16, 107.4, 106.6, 105.88, 105.16, 104.16, 103.36, 102.48, 101.52, 100.56, 99.72, 98.6, 97.68, 96.64, 95.68, 93.96, 92.76, 91.16, 89.92, 88.72, 87.52, 86.32, 84.96, 83.76, 82.08, 80.68, 79.44, 77.72, 76.36, 74.52, 73.24, 71.88, 70.28, 68.84, 67.68, 66.0, 64.64, 63.48, 62.0, 60.76, 59.72, 58.32, 57.24, 56.24, 55.0, 53.92, 53.04, 51.72, 50.6, 49.56, 48.4, 47.04, 45.76, 44.6, 43.0, 41.64, 40.52, 38.96, 37.6, 36.32, 34.68, 33.28, 32.16, 30.44, 29.16, 28.12, 26.64, 25.44, 24.44, 23.04, 21.88, 20.84, 19.48, 18.28, 17.2, 15.96, 14.48, 13.32, 12.2, 10.56, 9.44, 8.0, 6.64, 5.44, 4.44, 3.04, 1.88, 111.52, 111.24, 110.68, 110.12, 109.56, 108.84, 108.24, 107.44, 106.72, 106.0, 105.08, 104.2, 103.36, 102.32, 101.36, 100.36, 99.4, 97.36, 96.04, 94.28, 92.84, 91.68, 90.2, 89.08, 87.68, 85.84, 84.56, 83.32, 81.8, 80.44, 79.28, 77.8, 76.48, 75.32, 73.72, 72.28, 71.04, 69.16, 67.72, 65.76, 64.2, 62.92, 61.12, 59.72, 58.12, 56.76, 55.6, 54.16, 52.84, 51.68, 50.24, 49.0, 47.84, 46.28, 44.92, 43.72, 42.12, 40.8, 39.72, 38.24, 37.12, 35.96, 34.44, 33.28, 32.12, 30.6, 29.4, 28.12, 26.8, 25.28, 24.08, 22.56, 21.32, 20.24, 18.92, 17.76, 16.76, 15.52, 14.16, 12.92, 11.84, 10.16, 8.6, 7.4, 6.16, 5.0, 4.0, 2.68, 1.52, 109.28, 108.92, 108.28, 107.68, 106.88, 106.24, 105.4, 104.72, 103.96, 103.12, 102.24, 101.4, 100.52, 99.6, 98.56, 97.68, 96.56, 94.96, 93.88, 92.44, 91.36, 90.36, 89.24, 88.24, 87.08, 85.96, 84.68, 83.28, 82.04, 80.84, 79.36, 78.04, 76.88, 74.92, 73.52, 71.8, 70.44, 69.2, 67.56, 66.16, 64.96, 63.16, 61.8, 60.52, 58.96, 57.56, 56.32, 54.72, 53.28, 51.76, 50.44, 49.24, 47.72, 46.52, 45.48, 43.8, 42.68, 41.6, 40.24, 39.12, 38.12, 37.0, 35.72, 34.64, 33.72, 32.28, 31.12, 30.08, 29.08, 27.68, 26.56, 25.56, 24.28, 23.16, 22.2, 21.08, 19.88, 18.8, 17.84, 16.56, 15.44, 14.32, 13.32, 12.0, 10.88, 9.96, 7.48, 6.48, 5.4, 4.12, 3.08, 2.08, 1.04, 107.52, 107.2, 106.64, 105.76, 105.0, 104.32, 103.4, 102.52, 101.76, 100.76, 99.8, 98.84, 97.92, 96.8, 96.04, 94.96, 93.8, 92.24, 91.0, 89.36, 88.12, 87.08, 85.88, 84.8, 83.6, 82.4, 81.0, 79.76, 78.64, 77.16, 75.84, 74.8, 73.28, 72.12, 70.88, 69.52, 68.32, 67.24, 65.96, 64.56, 63.24, 62.04, 60.52, 59.24, 58.12, 56.52, 55.16, 53.92, 52.24, 50.88, 49.68, 48.0, 46.68, 45.16, 43.84, 42.72, 41.28, 40.08, 39.0, 37.6, 36.32, 35.28, 34.08, 32.76, 31.56, 30.48, 28.96, 27.76, 26.8, 25.44, 24.36, 23.48, 22.32, 20.92, 19.88, 18.96, 17.76, 16.72, 15.8, 14.72, 13.36, 12.32, 11.2, 10.12, 7.72, 6.6, 5.4, 4.36, 3.36, 2.28, 1.12, 156.04, 155.0, 153.68, 152.24, 150.76, 149.12, 147.2, 145.24, 142.92, 139.72, 136.76, 134.08, 131.04, 127.76, 124.64, 121.48, 118.24, 114.72, 111.48, 108.56, 105.48, 102.6, 99.44, 96.56, 93.6, 90.8, 87.6, 84.68, 81.68, 78.84, 75.88, 73.16, 70.4, 67.84, 65.32, 62.68, 60.12, 57.48, 54.64, 51.68, 49.0, 46.28, 43.84, 41.44, 38.84, 36.52, 33.92, 31.6, 29.16, 26.52, 24.0, 21.48, 18.96, 16.72, 14.04, 11.72, 9.16, 6.4, 4.16, 1.88, 163.8, 162.6, 161.32, 159.84, 158.44, 156.76, 154.88, 153.0, 150.6, 147.24, 143.96, 141.04, 137.64, 134.2, 130.84, 127.92, 124.92, 121.88, 119.04, 116.12, 113.04, 110.32, 107.44, 104.72, 101.8, 99.12, 96.4, 93.64, 91.08, 88.44, 85.76, 83.24, 80.52, 77.6, 74.8, 71.8, 68.72, 65.6, 62.8, 60.04, 57.16, 54.48, 51.52, 48.92, 46.28, 43.88, 41.52, 39.16, 37.0, 34.72, 32.68, 30.16, 27.76, 25.28, 22.84, 20.4, 17.92, 15.68, 13.32, 11.08, 8.52, 6.16, 4.0, 1.88, 150.44, 149.2, 147.76, 146.2, 144.56, 142.84, 141.12, 139.12, 136.64, 133.52, 130.76, 128.28, 125.76, 122.92, 120.08, 117.48, 114.88, 112.12, 109.56, 106.96, 104.2, 101.72, 99.08, 96.36, 93.36, 90.68, 87.88, 85.44, 82.88, 80.28, 78.0, 75.4, 72.92, 70.36, 67.64, 65.04, 62.32, 59.52, 56.92, 54.24, 51.52, 49.0, 46.64, 44.16, 41.8, 39.2, 36.76, 34.44, 32.08, 29.72, 27.48, 25.16, 22.72, 20.2, 17.88, 15.52, 13.08, 10.76, 7.28, 5.08, 2.8, 1.0, 183.08, 181.88, 180.48, 178.96, 177.32, 175.68, 173.84, 171.92, 169.6, 166.6, 163.84, 161.4, 159.0, 156.24, 153.8, 151.28, 148.72, 146.24, 143.68, 141.04, 138.48, 135.84, 133.2, 130.72, 128.2, 125.6, 123.12, 120.36, 117.88, 115.32, 112.6, 110.08, 107.48, 104.84, 102.36, 99.92, 97.28, 94.84, 92.48, 90.12, 87.8, 85.24, 82.88, 80.4, 77.88, 75.32, 72.68, 70.2, 67.56, 64.84, 62.28, 59.68, 57.08, 54.76, 52.4, 49.96, 47.52, 44.92, 42.52, 40.12, 37.72, 35.68, 33.44, 31.48, 29.04, 26.8, 24.52, 22.24, 19.92, 17.52, 15.44, 12.92, 10.68, 8.08, 5.84, 3.84, 2.0, 207.64, 206.56, 205.2, 203.76, 202.2, 200.56, 198.8, 196.96, 194.84, 192.08, 189.4, 187.0, 184.52, 181.72, 179.04, 176.24, 173.32, 170.24, 167.48, 164.6, 161.6, 158.88, 156.12, 153.36, 150.52, 147.84, 145.12, 142.32, 139.6, 136.76, 133.88, 131.24, 128.56, 125.84, 123.28, 120.72, 118.12, 115.68, 113.12, 110.44, 107.8, 105.04, 102.24, 99.6, 97.0, 94.24, 91.76, 89.32, 86.76, 84.56, 82.04, 79.72, 77.28, 74.68, 72.28, 69.32, 66.36, 63.76, 61.08, 58.4, 55.96, 53.44, 50.8, 48.56, 46.2, 43.92, 41.44, 38.76, 36.52, 33.84, 31.28, 28.84, 26.48, 24.16, 21.84, 19.4, 17.08, 14.64, 12.4, 9.96, 7.56, 5.4, 3.04, 1.56, 209.16, 207.92, 206.44, 204.84, 203.24, 201.52, 199.68, 197.64, 195.24, 192.44, 189.88, 187.68, 185.44, 182.88, 180.4, 177.88, 175.32, 172.64, 169.88, 167.32, 164.72, 161.96, 159.36, 156.68, 153.88, 151.32, 148.64, 145.8, 143.16, 140.2, 137.4, 134.56, 131.8, 128.92, 125.88, 123.12, 120.16, 117.36, 114.6, 112.04, 109.32, 106.52, 103.88, 101.16, 98.48, 96.04, 93.56, 90.92, 88.44, 85.76, 83.08, 80.64, 77.8, 75.0, 72.12, 69.4, 66.48, 63.72, 61.0, 58.2, 55.64, 53.12, 50.44, 48.04, 45.56, 42.96, 40.48, 37.88, 35.28, 32.68, 30.08, 27.8, 25.64, 23.36, 21.28, 18.88, 16.72, 14.52, 12.36, 9.92, 7.44, 5.2, 2.84, 1.32, 207.8, 206.56, 205.12, 203.56, 201.96, 200.16, 198.36, 196.32, 193.88, 191.12, 188.68, 186.44, 184.24, 181.68, 179.4, 176.68, 174.12, 171.48, 168.88, 166.36, 163.68, 161.2, 158.6, 155.88, 153.16, 150.68, 148.16, 145.48, 142.8, 140.16, 137.44, 135.0, 132.36, 129.68, 127.36, 124.76, 122.36, 119.8, 117.2, 114.8, 112.48, 110.24, 107.76, 105.24, 102.64, 99.92, 97.2, 94.68, 92.12, 89.44, 87.0, 84.56, 82.12, 79.72, 77.28, 75.0, 72.72, 70.32, 67.92, 65.36, 62.88, 60.24, 57.56, 55.08, 52.56, 50.04, 47.64, 45.2, 42.96, 40.64, 38.4, 36.04, 33.6, 31.32, 29.0, 26.72, 24.36, 21.8, 19.6, 17.12, 14.92, 12.6, 10.2, 7.64, 5.32, 3.24, 1.52, 296.08, 293.68, 290.72, 287.12, 282.0, 275.92, 270.08, 264.24, 258.64, 252.96, 247.28, 241.52, 235.76, 229.92, 224.0, 218.32, 212.4, 206.88, 201.36, 196.0, 190.4, 184.72, 178.88, 173.12, 167.52, 162.16, 156.96, 152.0, 146.88, 141.76, 136.56, 131.44, 126.16, 120.72, 114.88, 108.96, 103.36, 97.92, 93.04, 88.08, 83.12, 77.68, 72.56, 67.68, 62.64, 57.84, 53.28, 48.32, 43.36, 38.24, 33.28, 28.56, 24.0, 19.44, 14.8, 9.84, 5.2, 2.0, 312.32, 309.44, 306.08, 302.24, 297.28, 291.44, 285.76, 279.76, 273.68, 267.12, 260.4, 253.92, 247.92, 241.92, 236.16, 230.4, 224.64, 219.12, 213.6, 208.08, 202.52, 196.84, 191.4, 185.96, 180.68, 175.32, 169.64, 163.56, 157.96, 152.44, 147.16, 142.04, 137.0, 132.04, 127.16, 122.28, 117.24, 112.04, 106.92, 101.72, 96.8, 91.76, 86.48, 81.04, 75.92, 70.88, 65.44, 60.24, 55.6, 50.64, 45.6, 40.48, 35.04, 29.76, 24.64, 19.84, 14.96, 10.32, 5.44, 2.16, 334.88, 332.0, 328.88, 325.2, 320.4, 315.12, 310.24, 305.2, 299.92, 294.64, 289.28, 283.68, 278.24, 272.88, 267.28, 261.76, 256.24, 250.72, 245.36, 239.92, 234.68, 229.32, 223.88, 218.76, 213.72, 208.68, 203.72, 198.76, 193.72, 188.6, 183.4, 178.12, 172.84, 167.48, 162.28, 157.16, 152.12, 147.0, 142.2, 137.24, 132.2, 127.08, 122.12, 117.08, 112.04, 107.24, 102.76, 98.28, 93.64, 89.08, 84.44, 79.64, 74.52, 69.72, 64.76, 60.04, 55.48, 51.0, 46.52, 41.64, 36.68, 31.76, 27.16, 22.8, 18.36, 13.88, 9.16, 4.6, 1.92, 374.28, 371.96, 369.0, 365.4, 360.6, 355.48, 350.84, 345.96, 340.84, 335.96, 331.4, 326.68, 321.96, 317.32, 312.44, 307.24, 302.12, 296.92, 291.64, 286.28, 280.8, 275.2, 269.92, 264.64, 259.44, 254.32, 249.44, 244.4, 239.52, 234.64, 229.92, 225.36, 220.88, 216.4, 211.92, 207.04, 202.24, 197.28, 192.4, 187.52, 182.56, 177.68, 172.8, 167.76, 162.88, 157.92, 153.12, 148.16, 143.28, 138.24, 133.04, 127.92, 122.96, 118.0, 112.96, 107.84, 102.88, 98.24, 93.76, 89.04, 84.28, 79.8, 75.12, 70.56, 66.0, 61.4, 56.96, 52.68, 48.16, 43.52, 38.92, 34.6, 30.36, 26.16, 21.88, 17.52, 13.08, 8.6, 4.52, 1.88, 407.12, 404.56, 401.6, 398.24, 393.6, 388.8, 384.32, 379.28, 374.0, 368.8, 363.68, 358.72, 353.84, 349.04, 344.16, 339.12, 333.76, 328.56, 323.44, 318.24, 313.32, 308.36, 303.4, 298.44, 293.24, 288.2, 283.16, 278.2, 273.08, 267.96, 263.08, 258.12, 253.24, 248.52, 243.88, 239.32, 234.76, 230.12, 225.32, 220.68, 215.92, 211.2, 206.32, 201.44, 196.72, 192.08, 187.28, 182.48, 177.76, 172.96, 168.24, 163.6, 158.8, 154.16, 149.52, 144.88, 140.16, 135.44, 130.56, 125.44, 120.32, 115.2, 109.92, 104.88, 100.08, 95.2, 90.24, 85.2, 80.16, 75.36, 70.32, 65.28, 60.72, 56.16, 51.84, 47.12, 42.32, 37.6, 32.88, 28.48, 24.12, 19.8, 15.32, 10.84, 6.4, 2.72, 405.92, 403.04, 399.68, 395.84, 390.88, 385.68, 380.96, 376.16, 371.28, 366.56, 361.92, 357.28, 352.72, 348.0, 343.36, 338.56, 333.92, 329.12, 324.4, 319.76, 315.0, 310.12, 305.32, 300.44, 295.64, 290.68, 285.8, 280.68, 275.56, 270.36, 265.16, 260.04, 254.76, 249.72, 244.68, 239.64, 234.52, 229.4, 224.2, 219.08, 214.0, 208.88, 203.68, 198.56, 193.52, 188.64, 183.84, 178.96, 174.24, 169.6, 165.04, 160.4, 155.76, 151.04, 146.4, 141.92, 137.12, 132.64, 128.48, 124.0, 119.0, 114.12, 109.2, 104.28, 99.32, 94.56, 90.16, 85.68, 81.28, 76.88, 72.36, 68.08, 63.72, 59.4, 55.2, 50.88, 46.72, 42.48, 37.92, 33.36, 29.04, 24.56, 20.32, 16.08, 12.0, 6.64, 2.56, 506.08, 502.0, 496.96, 489.84, 482.72, 475.04, 467.2, 459.44, 451.68, 444.0, 436.32, 428.56, 420.32, 412.32, 404.48, 396.56, 388.56, 380.64, 372.72, 364.96, 357.04, 349.12, 341.44, 333.92, 326.64, 319.44, 312.16, 305.04, 297.84, 290.48, 283.12, 275.84, 268.64, 261.36, 254.16, 246.64, 239.36, 232.0, 224.72, 217.68, 210.76, 203.8, 196.76, 189.72, 182.52, 175.48, 168.36, 161.48, 154.68, 147.72, 140.68, 133.96, 126.92, 119.72, 112.44, 105.0, 97.72, 90.52, 83.32, 76.2, 68.96, 62.0, 55.36, 48.88, 42.48, 36.32, 30.0, 23.68, 18.08, 12.32, 6.56, 2.08}
    pres_qc = 
      {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
    psal = 
      {34.0, 34.0, 34.0, 34.0, 34.0, 33.872, 33.856, 33.848, 33.849, 33.844, 33.839, 33.831, 33.829, 33.826, 33.825, 33.824, 33.822, 33.822, 33.815, 33.807, 33.805, 33.79, 33.783, 33.767, 33.755, 33.75, 33.742, 33.74, 33.735, 33.731, 33.728, 33.723, 33.706, 33.644, 33.593, 33.562, 33.547, 33.518, 33.509, 33.502, 33.478, 33.454, 33.44, 33.441, 33.441, 33.44, 33.439, 33.437, 33.427, 33.414, 33.401, 33.346, 33.335, 33.326, 33.308, 33.245, 33.225, 33.192, 33.121, 33.06, 32.996, 32.94, 32.936, 32.899, 32.879, 32.828, 32.784, 32.773, 32.767, 32.76, 32.756, 32.753, 32.752, 32.751, 32.751, 32.751, 32.749, 32.747, 32.743, 32.723, 32.71, 32.699, 32.696, 32.683, 32.652, 32.648, 32.638, 32.636, 32.631, 32.629, 32.623, 32.618, 32.614, 32.597, 32.594, 32.593, 32.596, 32.589, 32.574, 32.55, 32.555, 33.847, 33.847, 33.847, 33.846, 33.845, 33.846, 33.844, 33.844, 33.842, 33.837, 33.824, 33.815, 33.789, 33.774, 33.768, 33.761, 33.757, 33.753, 33.752, 33.741, 33.7, 33.683, 33.651, 33.652, 33.631, 33.625, 33.618, 33.605, 33.588, 33.572, 33.564, 33.555, 33.552, 33.548, 33.536, 33.512, 33.509, 33.509, 33.503, 33.478, 33.453, 33.44, 33.428, 33.427, 33.404, 33.397, 33.331, 33.269, 33.263, 33.214, 33.141, 33.064, 33.023, 32.962, 32.939, 32.934, 32.932, 32.931, 32.905, 32.867, 32.818, 32.785, 32.774, 32.769, 32.767, 32.764, 32.76, 32.753, 32.741, 32.729, 32.712, 32.695, 32.691, 32.678, 32.645, 32.606, 32.574, 32.558, 32.56, 32.56, 32.56, 32.56, 32.558, 32.559, 32.558, 32.558, 32.556, 32.558, 32.557, 33.855, 33.855, 33.854, 33.849, 33.834, 33.823, 33.82, 33.803, 33.785, 33.775, 33.767, 33.763, 33.761, 33.755, 33.755, 33.755, 33.757, 33.758, 33.757, 33.746, 33.724, 33.706, 33.667, 33.651, 33.634, 33.617, 33.613, 33.608, 33.603, 33.602, 33.598, 33.593, 33.579, 33.555, 33.535, 33.524, 33.505, 33.491, 33.451, 33.431, 33.434, 33.433, 33.423, 33.4, 33.379, 33.338, 33.258, 33.211, 33.164, 33.135, 33.12, 33.112, 33.109, 33.109, 33.109, 33.11, 33.107, 33.045, 32.985, 32.939, 32.938, 32.94, 32.94, 32.89, 32.872, 32.831, 32.784, 32.768, 32.759, 32.753, 32.742, 32.726, 32.713, 32.698, 32.644, 32.592, 32.568, 32.554, 32.551, 32.55, 32.551, 32.548, 32.548, 32.547, 32.546, 32.547, 32.548, 32.545, 32.546, 33.806, 33.803, 33.787, 33.774, 33.758, 33.752, 33.751, 33.75, 33.747, 33.728, 33.711, 33.701, 33.693, 33.681, 33.672, 33.669, 33.667, 33.655, 33.646, 33.633, 33.623, 33.61, 33.6, 33.599, 33.587, 33.583, 33.577, 33.574, 33.57, 33.569, 33.556, 33.547, 33.541, 33.535, 33.529, 33.519, 33.508, 33.501, 33.472, 33.458, 33.444, 33.409, 33.359, 33.289, 33.256, 33.237, 33.196, 33.164, 33.144, 33.131, 33.122, 33.103, 33.075, 33.043, 33.044, 33.017, 33.003, 33.003, 32.981, 32.968, 32.95, 32.915, 32.904, 32.871, 32.846, 32.828, 32.819, 32.812, 32.805, 32.788, 32.782, 32.778, 32.766, 32.753, 32.732, 32.72, 32.679, 32.632, 32.581, 32.559, 32.555, 32.549, 32.549, 32.55, 32.549, 32.549, 32.55, 32.549, 32.549, 32.546, 32.546, 32.546, 32.544, 33.769, 33.769, 33.759, 33.746, 33.735, 33.727, 33.724, 33.718, 33.718, 33.711, 33.709, 33.704, 33.703, 33.701, 33.695, 33.683, 33.681, 33.673, 33.666, 33.66, 33.656, 33.655, 33.648, 33.646, 33.644, 33.64, 33.631, 33.629, 33.627, 33.612, 33.598, 33.567, 33.536, 33.528, 33.521, 33.5, 33.484, 33.486, 33.437, 33.423, 33.417, 33.39, 33.327, 33.274, 33.203, 33.172, 33.12, 33.11, 33.104, 33.104, 33.107, 33.073, 33.048, 32.989, 32.972, 32.957, 32.943, 32.907, 32.888, 32.851, 32.836, 32.834, 32.824, 32.831, 32.821, 32.813, 32.801, 32.779, 32.77, 32.754, 32.719, 32.709, 32.698, 32.656, 32.599, 32.578, 32.562, 32.551, 32.551, 32.55, 32.551, 32.551, 32.552, 32.554, 32.552, 32.552, 32.55, 32.55, 32.549, 32.549, 32.54, 33.916, 33.917, 33.918, 33.918, 33.92, 33.919, 33.918, 33.917, 33.917, 33.917, 33.915, 33.896, 33.88, 33.877, 33.877, 33.855, 33.847, 33.846, 33.839, 33.838, 33.837, 33.833, 33.828, 33.818, 33.795, 33.74, 33.708, 33.694, 33.678, 33.673, 33.666, 33.658, 33.633, 33.529, 33.514, 33.509, 33.485, 33.412, 33.293, 33.255, 33.202, 33.156, 33.096, 33.032, 32.89, 32.854, 32.838, 32.78, 32.704, 32.666, 32.632, 32.6, 32.576, 32.568, 32.556, 32.554, 32.558, 32.56, 32.554, 32.546, 33.934, 33.935, 33.935, 33.936, 33.936, 33.935, 33.935, 33.934, 33.936, 33.929, 33.926, 33.926, 33.927, 33.927, 33.928, 33.928, 33.916, 33.911, 33.891, 33.878, 33.879, 33.872, 33.864, 33.857, 33.849, 33.848, 33.824, 33.786, 33.749, 33.733, 33.694, 33.685, 33.677, 33.67, 33.655, 33.556, 33.509, 33.497, 33.496, 33.492, 33.472, 33.45, 33.376, 33.32, 33.296, 33.19, 33.06, 32.992, 32.894, 32.848, 32.752, 32.662, 32.614, 32.606, 32.598, 32.592, 32.582, 32.57, 32.564, 32.564, 32.564, 32.564, 32.564, 32.554, 33.949, 33.949, 33.95, 33.95, 33.95, 33.948, 33.947, 33.944, 33.941, 33.935, 33.936, 33.928, 33.916, 33.903, 33.903, 33.898, 33.89, 33.883, 33.867, 33.861, 33.862, 33.862, 33.842, 33.827, 33.822, 33.806, 33.779, 33.766, 33.746, 33.719, 33.703, 33.691, 33.683, 33.677, 33.632, 33.56, 33.541, 33.528, 33.519, 33.495, 33.422, 33.372, 33.346, 33.204, 33.072, 32.984, 32.964, 32.924, 32.902, 32.88, 32.79, 32.624, 32.584, 32.58, 32.584, 32.58, 32.574, 32.57, 32.564, 32.566, 32.557, 32.56, 34.023, 34.021, 34.02, 34.021, 34.02, 34.016, 34.013, 34.011, 34.008, 34.007, 34.006, 34.005, 34.003, 34.0, 33.996, 33.994, 33.987, 33.982, 33.98, 33.974, 33.964, 33.952, 33.936, 33.929, 33.923, 33.903, 33.892, 33.891, 33.89, 33.888, 33.886, 33.884, 33.874, 33.87, 33.867, 33.866, 33.848, 33.809, 33.781, 33.751, 33.729, 33.717, 33.705, 33.701, 33.695, 33.691, 33.685, 33.635, 33.557, 33.519, 33.511, 33.493, 33.449, 33.391, 33.341, 33.267, 33.097, 33.021, 33.019, 32.995, 32.936, 32.888, 32.854, 32.68, 32.568, 32.56, 32.564, 32.566, 32.566, 32.568, 32.566, 32.568, 32.566, 32.562, 32.564, 32.562, 32.562, 34.065, 34.065, 34.065, 34.065, 34.065, 34.065, 34.063, 34.06, 34.054, 34.04, 34.027, 34.02, 34.016, 34.014, 34.012, 34.008, 34.008, 34.01, 34.009, 34.006, 33.995, 33.991, 33.989, 33.979, 33.971, 33.97, 33.962, 33.954, 33.946, 33.939, 33.937, 33.92, 33.907, 33.903, 33.899, 33.897, 33.888, 33.877, 33.87, 33.865, 33.852, 33.845, 33.843, 33.84, 33.829, 33.79, 33.784, 33.776, 33.77, 33.759, 33.738, 33.71, 33.695, 33.643, 33.603, 33.573, 33.542, 33.521, 33.482, 33.435, 33.373, 33.287, 33.241, 33.221, 33.109, 33.083, 32.999, 32.859, 32.841, 32.795, 32.699, 32.627, 32.601, 32.599, 32.607, 32.617, 32.613, 32.607, 32.599, 32.591, 32.581, 32.575, 32.575, 32.576, 34.057, 34.057, 34.054, 34.05, 34.05, 34.047, 34.041, 34.033, 34.025, 34.019, 34.018, 34.016, 34.015, 34.016, 34.014, 34.015, 34.006, 33.997, 33.988, 33.985, 33.977, 33.974, 33.97, 33.97, 33.968, 33.967, 33.967, 33.967, 33.96, 33.922, 33.915, 33.912, 33.909, 33.91, 33.909, 33.904, 33.888, 33.887, 33.877, 33.872, 33.864, 33.851, 33.838, 33.828, 33.802, 33.791, 33.781, 33.773, 33.757, 33.715, 33.655, 33.621, 33.593, 33.566, 33.554, 33.546, 33.505, 33.468, 33.459, 33.42, 33.382, 33.334, 33.248, 33.216, 33.168, 33.112, 33.098, 33.094, 33.062, 32.966, 32.854, 32.726, 32.652, 32.606, 32.61, 32.608, 32.602, 32.598, 32.594, 32.59, 32.586, 32.574, 32.576, 32.576, 34.043, 34.038, 34.036, 34.035, 34.031, 34.025, 34.023, 34.021, 34.016, 34.012, 34.012, 34.006, 34.002, 34.002, 33.993, 33.988, 33.981, 33.978, 33.978, 33.978, 33.975, 33.975, 33.974, 33.965, 33.957, 33.954, 33.956, 33.956, 33.955, 33.953, 33.952, 33.935, 33.93, 33.923, 33.916, 33.914, 33.91, 33.904, 33.89, 33.882, 33.877, 33.874, 33.871, 33.86, 33.846, 33.844, 33.815, 33.8, 33.796, 33.79, 33.784, 33.782, 33.78, 33.769, 33.651, 33.608, 33.589, 33.564, 33.552, 33.513, 33.481, 33.449, 33.377, 33.233, 33.161, 33.137, 33.123, 33.109, 33.073, 33.059, 33.019, 32.857, 32.767, 32.753, 32.693, 32.659, 32.629, 32.613, 32.607, 32.597, 32.582, 32.576, 32.573, 32.572, 32.573, 32.573, 32.573, 34.099, 34.096, 34.09, 34.09, 34.087, 34.088, 34.084, 34.083, 34.079, 34.074, 34.074, 34.071, 34.07, 34.068, 34.064, 34.063, 34.041, 34.033, 34.027, 34.015, 34.008, 33.995, 33.988, 33.985, 33.977, 33.961, 33.952, 33.946, 33.937, 33.93, 33.915, 33.904, 33.884, 33.872, 33.856, 33.835, 33.811, 33.792, 33.78, 33.754, 33.6, 33.518, 33.468, 33.376, 33.18, 33.092, 33.078, 33.012, 32.978, 32.896, 32.81, 32.696, 32.63, 32.574, 32.568, 32.57, 32.57, 32.572, 34.106, 34.105, 34.102, 34.098, 34.096, 34.094, 34.091, 34.092, 34.093, 34.093, 34.091, 34.089, 34.079, 34.068, 34.065, 34.065, 34.059, 34.055, 34.041, 34.036, 34.028, 34.022, 34.017, 34.012, 34.004, 33.995, 33.986, 33.982, 33.974, 33.961, 33.949, 33.94, 33.929, 33.911, 33.895, 33.885, 33.864, 33.833, 33.8, 33.776, 33.756, 33.662, 33.56, 33.496, 33.45, 33.346, 33.26, 33.078, 33.074, 33.02, 32.956, 32.94, 32.908, 32.836, 32.692, 32.616, 32.574, 32.55, 32.538, 32.54, 34.109, 34.108, 34.109, 34.102, 34.099, 34.101, 34.1, 34.098, 34.098, 34.096, 34.096, 34.091, 34.093, 34.089, 34.083, 34.08, 34.072, 34.063, 34.061, 34.062, 34.058, 34.052, 34.046, 34.042, 34.038, 34.035, 34.02, 34.014, 34.012, 34.004, 33.987, 33.984, 33.974, 33.967, 33.96, 33.955, 33.939, 33.928, 33.894, 33.886, 33.858, 33.832, 33.828, 33.806, 33.794, 33.776, 33.766, 33.75, 33.668, 33.62, 33.536, 33.42, 33.318, 33.19, 33.122, 33.072, 32.978, 32.908, 32.804, 32.674, 32.6, 32.575, 32.572, 32.564, 32.559, 32.554, 32.554, 32.555, 32.555, 34.119, 34.121, 34.121, 34.121, 34.12, 34.118, 34.12, 34.118, 34.119, 34.115, 34.11, 34.11, 34.111, 34.111, 34.11, 34.108, 34.104, 34.103, 34.1, 34.09, 34.09, 34.092, 34.092, 34.088, 34.084, 34.08, 34.069, 34.069, 34.067, 34.061, 34.059, 34.055, 34.053, 34.047, 34.037, 34.039, 34.035, 34.018, 34.011, 34.001, 33.995, 33.977, 33.967, 33.962, 33.956, 33.947, 33.924, 33.906, 33.899, 33.857, 33.848, 33.842, 33.834, 33.818, 33.78, 33.745, 33.728, 33.688, 33.596, 33.473, 33.389, 33.326, 33.23, 33.21, 33.189, 33.083, 32.983, 32.877, 32.839, 32.808, 32.744, 32.641, 32.602, 32.6, 32.598, 32.593, 32.59, 32.59, 32.583, 32.584, 34.135, 34.137, 34.137, 34.136, 34.136, 34.136, 34.134, 34.129, 34.126, 34.128, 34.126, 34.124, 34.121, 34.123, 34.122, 34.114, 34.113, 34.111, 34.107, 34.107, 34.103, 34.103, 34.101, 34.101, 34.098, 34.098, 34.095, 34.088, 34.082, 34.077, 34.072, 34.07, 34.062, 34.057, 34.05, 34.047, 34.047, 34.042, 34.039, 34.032, 34.027, 34.025, 34.016, 34.012, 34.004, 33.998, 33.993, 33.979, 33.958, 33.959, 33.952, 33.953, 33.94, 33.917, 33.908, 33.891, 33.878, 33.86, 33.835, 33.804, 33.78, 33.762, 33.729, 33.711, 33.696, 33.66, 33.585, 33.579, 33.561, 33.522, 33.483, 33.438, 33.36, 33.264, 33.006, 32.808, 32.781, 32.76, 32.751, 32.763, 32.755, 32.673, 32.665, 32.637, 32.631, 32.632, 34.134, 34.134, 34.132, 34.127, 34.128, 34.127, 34.125, 34.123, 34.122, 34.121, 34.12, 34.12, 34.119, 34.118, 34.114, 34.11, 34.108, 34.106, 34.105, 34.104, 34.101, 34.101, 34.101, 34.097, 34.092, 34.09, 34.088, 34.084, 34.083, 34.079, 34.073, 34.071, 34.065, 34.055, 34.045, 34.036, 34.031, 34.023, 34.021, 34.025, 34.028, 34.028, 34.02, 34.015, 34.004, 33.993, 33.982, 33.982, 33.976, 33.968, 33.959, 33.943, 33.912, 33.894, 33.87, 33.852, 33.853, 33.854, 33.84, 33.811, 33.8, 33.798, 33.792, 33.744, 33.694, 33.664, 33.644, 33.65, 33.622, 33.51, 33.474, 33.362, 33.306, 33.226, 33.14, 33.016, 32.884, 32.762, 32.712, 32.65, 32.613, 32.59, 32.57, 32.569, 32.571, 32.574, 32.574, 34.174, 34.174, 34.17, 34.166, 34.16, 34.159, 34.156, 34.148, 34.144, 34.136, 34.132, 34.133, 34.134, 34.134, 34.128, 34.123, 34.123, 34.121, 34.117, 34.118, 34.117, 34.117, 34.114, 34.108, 34.1, 34.1, 34.1, 34.102, 34.103, 34.095, 34.091, 34.072, 34.062, 34.054, 34.033, 34.03, 34.026, 34.016, 34.011, 34.007, 34.007, 34.006, 34.001, 33.99, 33.982, 33.974, 33.973, 33.946, 33.911, 33.896, 33.877, 33.866, 33.834, 33.805, 33.79, 33.777, 33.766, 33.743, 33.68, 33.604, 33.558, 33.386, 33.216, 32.992, 32.874, 32.796, 32.796, 32.668, 32.548, 32.52, 32.528, 32.53}
    psal_qc = 
      {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
    temp = 
      {10.133, 11.679, 12.906, 14.508, 15.446, 9.502, 9.564, 9.614, 9.628, 9.662, 9.695, 9.71, 9.719, 9.725, 9.729, 9.733, 9.739, 9.74, 9.756, 9.765, 9.769, 9.793, 9.796, 9.809, 9.82, 9.822, 9.818, 9.82, 9.824, 9.839, 9.846, 9.854, 9.836, 9.765, 9.713, 9.763, 9.769, 9.837, 9.895, 9.93, 9.999, 10.102, 10.17, 10.186, 10.198, 10.225, 10.255, 10.282, 10.336, 10.39, 10.417, 10.498, 10.501, 10.516, 10.537, 10.558, 10.588, 10.555, 10.414, 10.321, 10.39, 10.312, 10.621, 10.852, 10.951, 10.944, 10.909, 10.908, 10.909, 10.9, 10.892, 10.888, 10.887, 10.886, 10.886, 10.886, 10.888, 10.889, 10.883, 10.876, 10.885, 10.902, 10.915, 10.948, 11.013, 11.025, 11.06, 11.07, 11.082, 11.088, 11.106, 11.126, 11.143, 11.187, 11.196, 11.194, 11.191, 11.212, 11.275, 11.304, 11.287, 9.647, 9.65, 9.653, 9.658, 9.663, 9.666, 9.669, 9.675, 9.685, 9.705, 9.737, 9.761, 9.79, 9.804, 9.811, 9.834, 9.861, 9.893, 9.908, 9.905, 9.84, 9.798, 9.727, 9.73, 9.716, 9.718, 9.729, 9.73, 9.734, 9.755, 9.768, 9.788, 9.793, 9.804, 9.836, 9.904, 9.916, 9.925, 9.942, 10.03, 10.134, 10.23, 10.323, 10.362, 10.425, 10.443, 10.467, 10.446, 10.446, 10.446, 10.317, 10.236, 10.248, 10.257, 10.26, 10.356, 10.632, 10.755, 10.872, 10.914, 10.917, 10.903, 10.898, 10.89, 10.884, 10.881, 10.885, 10.872, 10.868, 10.87, 10.893, 10.935, 10.948, 10.977, 11.069, 11.17, 11.262, 11.312, 11.314, 11.326, 11.332, 11.339, 11.354, 11.358, 11.39, 11.379, 11.399, 11.402, 11.411, 9.623, 9.625, 9.629, 9.647, 9.703, 9.735, 9.744, 9.771, 9.796, 9.806, 9.817, 9.827, 9.833, 9.845, 9.854, 9.862, 9.87, 9.898, 9.912, 9.893, 9.837, 9.797, 9.735, 9.709, 9.699, 9.701, 9.703, 9.703, 9.701, 9.699, 9.697, 9.703, 9.719, 9.767, 9.833, 9.859, 9.921, 9.971, 10.131, 10.315, 10.33, 10.356, 10.405, 10.453, 10.473, 10.475, 10.419, 10.364, 10.305, 10.27, 10.265, 10.258, 10.256, 10.252, 10.252, 10.251, 10.247, 10.216, 10.186, 10.24, 10.24, 10.246, 10.513, 10.729, 10.843, 10.891, 10.897, 10.873, 10.873, 10.861, 10.861, 10.882, 10.906, 10.936, 11.074, 11.206, 11.254, 11.293, 11.308, 11.335, 11.346, 11.369, 11.371, 11.388, 11.408, 11.418, 11.43, 11.454, 11.465, 9.791, 9.794, 9.805, 9.811, 9.817, 9.868, 9.88, 9.898, 9.905, 9.87, 9.816, 9.784, 9.762, 9.744, 9.732, 9.723, 9.721, 9.705, 9.693, 9.689, 9.693, 9.707, 9.721, 9.729, 9.775, 9.789, 9.809, 9.819, 9.835, 9.843, 9.879, 9.903, 9.917, 9.915, 9.919, 9.943, 9.965, 9.989, 10.113, 10.267, 10.368, 10.432, 10.444, 10.424, 10.38, 10.364, 10.32, 10.292, 10.324, 10.352, 10.368, 10.464, 10.448, 10.376, 10.412, 10.84, 10.796, 10.792, 10.808, 10.808, 10.823, 10.889, 10.912, 10.917, 10.908, 10.903, 10.9, 10.897, 10.896, 10.883, 10.876, 10.872, 10.865, 10.86, 10.879, 10.902, 10.999, 11.11, 11.226, 11.293, 11.304, 11.309, 11.318, 11.321, 11.337, 11.342, 11.366, 11.374, 11.406, 11.437, 11.444, 11.461, 11.517, 9.78, 9.78, 9.792, 9.809, 9.809, 9.813, 9.813, 9.808, 9.808, 9.802, 9.799, 9.784, 9.785, 9.777, 9.773, 9.753, 9.736, 9.728, 9.721, 9.72, 9.722, 9.72, 9.724, 9.726, 9.728, 9.73, 9.734, 9.738, 9.74, 9.76, 9.796, 9.906, 10.002, 10.032, 10.056, 10.106, 10.154, 10.218, 10.398, 10.418, 10.426, 10.444, 10.438, 10.384, 10.34, 10.382, 10.582, 10.62, 10.67, 10.69, 10.71, 10.862, 10.862, 10.864, 10.86, 10.858, 10.866, 10.876, 10.872, 10.866, 10.865, 10.865, 10.865, 10.864, 10.863, 10.864, 10.864, 10.867, 10.871, 10.877, 10.907, 10.924, 10.975, 11.073, 11.195, 11.246, 11.289, 11.331, 11.342, 11.346, 11.348, 11.355, 11.362, 11.379, 11.417, 11.43, 11.447, 11.459, 11.468, 11.531, 11.634, 9.072, 9.074, 9.074, 9.074, 9.074, 9.072, 9.074, 9.072, 9.072, 9.074, 9.078, 9.22, 9.368, 9.424, 9.428, 9.548, 9.6, 9.61, 9.644, 9.662, 9.667, 9.685, 9.706, 9.724, 9.736, 9.736, 9.718, 9.715, 9.709, 9.712, 9.715, 9.724, 9.766, 10.09, 10.147, 10.165, 10.255, 10.402, 10.381, 10.342, 10.348, 10.45, 10.807, 10.84, 10.834, 10.843, 10.849, 10.861, 10.963, 11.05, 11.167, 11.221, 11.269, 11.308, 11.332, 11.344, 11.383, 11.431, 11.515, 11.632, 8.919, 8.919, 8.921, 8.919, 8.923, 8.923, 8.927, 8.923, 8.937, 8.971, 8.983, 8.989, 8.985, 8.983, 8.979, 8.989, 9.079, 9.121, 9.293, 9.423, 9.451, 9.489, 9.527, 9.577, 9.619, 9.637, 9.709, 9.729, 9.719, 9.719, 9.705, 9.711, 9.715, 9.719, 9.741, 9.987, 10.187, 10.255, 10.263, 10.271, 10.309, 10.345, 10.384, 10.375, 10.366, 10.276, 10.597, 10.771, 10.783, 10.837, 10.987, 11.197, 11.284, 11.299, 11.296, 11.296, 11.302, 11.326, 11.338, 11.35, 11.418, 11.442, 11.494, 11.648, 8.834, 8.836, 8.836, 8.839, 8.841, 8.851, 8.852, 8.869, 8.894, 8.926, 8.95, 8.997, 9.103, 9.208, 9.244, 9.295, 9.36, 9.41, 9.497, 9.539, 9.545, 9.557, 9.645, 9.689, 9.699, 9.713, 9.731, 9.727, 9.729, 9.727, 9.725, 9.721, 9.721, 9.723, 9.799, 9.951, 10.051, 10.123, 10.167, 10.225, 10.318, 10.369, 10.372, 10.27, 10.327, 10.579, 10.684, 10.699, 10.744, 10.798, 10.948, 11.281, 11.386, 11.401, 11.401, 11.407, 11.413, 11.422, 11.437, 11.479, 11.626, 11.635, 8.333, 8.362, 8.374, 8.382, 8.394, 8.419, 8.435, 8.442, 8.462, 8.48, 8.495, 8.51, 8.529, 8.564, 8.587, 8.608, 8.66, 8.688, 8.71, 8.75, 8.798, 8.866, 8.944, 8.98, 9.026, 9.208, 9.29, 9.342, 9.368, 9.394, 9.422, 9.446, 9.508, 9.536, 9.552, 9.564, 9.608, 9.674, 9.71, 9.724, 9.735, 9.737, 9.733, 9.731, 9.729, 9.727, 9.727, 9.793, 9.945, 10.103, 10.137, 10.191, 10.259, 10.325, 10.353, 10.297, 10.165, 10.233, 10.363, 10.611, 10.614, 10.725, 10.824, 11.133, 11.46, 11.502, 11.514, 11.532, 11.55, 11.559, 11.559, 11.565, 11.58, 11.655, 11.697, 11.709, 11.712, 7.957, 7.961, 7.975, 7.984, 7.987, 7.989, 7.991, 8.008, 8.058, 8.173, 8.263, 8.327, 8.37, 8.401, 8.436, 8.472, 8.485, 8.487, 8.502, 8.529, 8.616, 8.654, 8.662, 8.698, 8.724, 8.742, 8.78, 8.812, 8.844, 8.888, 8.914, 9.05, 9.194, 9.258, 9.32, 9.37, 9.446, 9.496, 9.526, 9.552, 9.593, 9.613, 9.621, 9.629, 9.651, 9.727, 9.735, 9.737, 9.739, 9.735, 9.755, 9.763, 9.761, 9.731, 9.729, 9.777, 9.955, 10.087, 10.205, 10.279, 10.288, 10.234, 10.183, 10.174, 10.159, 10.381, 10.651, 10.852, 10.876, 10.957, 11.107, 11.341, 11.47, 11.548, 11.587, 11.644, 11.692, 11.707, 11.725, 11.749, 11.787, 11.802, 11.806, 11.808, 8.07, 8.081, 8.123, 8.159, 8.168, 8.182, 8.211, 8.258, 8.311, 8.363, 8.385, 8.409, 8.416, 8.428, 8.442, 8.465, 8.538, 8.617, 8.688, 8.735, 8.795, 8.829, 8.857, 8.867, 8.867, 8.865, 8.869, 8.879, 8.893, 9.089, 9.173, 9.241, 9.285, 9.299, 9.311, 9.357, 9.457, 9.471, 9.503, 9.523, 9.555, 9.601, 9.645, 9.679, 9.737, 9.755, 9.779, 9.797, 9.795, 9.727, 9.559, 9.539, 9.591, 9.755, 9.873, 9.939, 10.129, 10.259, 10.281, 10.287, 10.277, 10.249, 10.157, 10.121, 10.081, 10.125, 10.205, 10.285, 10.709, 10.821, 10.917, 11.061, 11.313, 11.533, 11.573, 11.589, 11.597, 11.589, 11.577, 11.561, 11.55, 11.652, 11.675, 11.669, 8.225, 8.286, 8.334, 8.351, 8.399, 8.435, 8.442, 8.446, 8.47, 8.509, 8.524, 8.57, 8.595, 8.608, 8.656, 8.703, 8.77, 8.819, 8.835, 8.842, 8.881, 8.877, 8.906, 8.957, 9.045, 9.076, 9.079, 9.086, 9.1, 9.12, 9.128, 9.211, 9.25, 9.285, 9.31, 9.323, 9.341, 9.375, 9.453, 9.486, 9.505, 9.517, 9.529, 9.565, 9.61, 9.622, 9.7, 9.745, 9.76, 9.778, 9.793, 9.802, 9.811, 9.823, 9.622, 9.553, 9.574, 9.673, 9.814, 10.132, 10.262, 10.266, 10.254, 10.082, 9.97, 9.998, 10.134, 10.234, 10.326, 10.546, 10.618, 11.042, 11.042, 11.082, 11.206, 11.306, 11.43, 11.506, 11.538, 11.554, 11.571, 11.6, 11.639, 11.654, 11.659, 11.662, 11.657, 7.425, 7.495, 7.577, 7.597, 7.631, 7.667, 7.731, 7.771, 7.819, 7.891, 7.911, 7.953, 7.985, 8.017, 8.051, 8.067, 8.197, 8.285, 8.329, 8.433, 8.483, 8.595, 8.681, 8.729, 8.807, 9.003, 9.121, 9.175, 9.225, 9.259, 9.311, 9.357, 9.449, 9.497, 9.581, 9.657, 9.735, 9.787, 9.825, 9.863, 9.66, 9.836, 9.984, 9.972, 9.944, 10.364, 10.612, 10.5, 10.86, 11.02, 11.14, 11.392, 11.488, 11.54, 11.592, 11.62, 11.632, 11.632, 7.295, 7.329, 7.381, 7.425, 7.459, 7.495, 7.543, 7.555, 7.553, 7.561, 7.589, 7.633, 7.779, 7.943, 8.015, 8.031, 8.113, 8.159, 8.251, 8.287, 8.343, 8.385, 8.427, 8.457, 8.493, 8.569, 8.667, 8.743, 8.871, 9.049, 9.141, 9.193, 9.253, 9.323, 9.391, 9.435, 9.523, 9.655, 9.781, 9.857, 9.897, 9.945, 9.853, 9.913, 9.965, 9.917, 9.825, 10.269, 10.569, 10.593, 10.673, 10.885, 10.953, 11.077, 11.397, 11.545, 11.613, 11.621, 11.621, 11.613, 7.186, 7.23, 7.232, 7.296, 7.354, 7.358, 7.368, 7.396, 7.41, 7.442, 7.47, 7.548, 7.57, 7.618, 7.704, 7.776, 7.878, 8.028, 8.13, 8.15, 8.204, 8.278, 8.328, 8.348, 8.378, 8.396, 8.462, 8.51, 8.532, 8.572, 8.722, 8.804, 8.936, 9.062, 9.132, 9.174, 9.198, 9.23, 9.336, 9.38, 9.521, 9.647, 9.675, 9.743, 9.791, 9.887, 9.931, 9.971, 10.087, 10.065, 10.021, 10.053, 10.127, 10.347, 10.511, 10.639, 10.875, 10.869, 11.051, 11.167, 11.356, 11.454, 11.472, 11.498, 11.562, 11.634, 11.641, 11.636, 11.631, 7.034, 7.034, 7.024, 7.032, 7.088, 7.135, 7.163, 7.219, 7.267, 7.316, 7.366, 7.373, 7.372, 7.374, 7.379, 7.394, 7.415, 7.435, 7.468, 7.582, 7.622, 7.64, 7.687, 7.751, 7.812, 7.856, 7.951, 7.98, 8.005, 8.047, 8.069, 8.122, 8.199, 8.25, 8.291, 8.346, 8.376, 8.396, 8.483, 8.559, 8.606, 8.738, 8.896, 9.074, 9.134, 9.166, 9.23, 9.292, 9.328, 9.508, 9.562, 9.582, 9.602, 9.65, 9.81, 10.004, 10.054, 10.112, 10.106, 10.034, 10.087, 10.201, 10.321, 10.387, 10.501, 10.666, 10.573, 10.51, 10.879, 11.119, 11.158, 11.377, 11.449, 11.443, 11.458, 11.479, 11.497, 11.518, 11.596, 11.602, 6.773, 6.771, 6.772, 6.77, 6.765, 6.773, 6.796, 6.857, 6.923, 6.94, 6.97, 7.015, 7.089, 7.119, 7.159, 7.19, 7.204, 7.238, 7.278, 7.302, 7.34, 7.422, 7.564, 7.618, 7.692, 7.754, 7.798, 7.842, 7.892, 7.94, 7.956, 7.984, 8.036, 8.098, 8.16, 8.18, 8.188, 8.206, 8.228, 8.298, 8.351, 8.357, 8.395, 8.429, 8.499, 8.579, 8.637, 8.741, 8.893, 9.007, 9.155, 9.183, 9.221, 9.259, 9.279, 9.335, 9.383, 9.415, 9.549, 9.677, 9.774, 9.826, 10.01, 10.162, 10.23, 10.286, 10.41, 10.458, 10.462, 10.422, 10.39, 10.374, 10.35, 10.334, 10.326, 9.874, 9.914, 10.358, 10.586, 10.882, 11.035, 11.261, 11.285, 11.381, 11.429, 11.431, 6.83, 6.843, 6.888, 6.933, 6.937, 6.954, 6.983, 7.032, 7.067, 7.085, 7.109, 7.116, 7.135, 7.164, 7.194, 7.239, 7.271, 7.3, 7.325, 7.347, 7.405, 7.435, 7.489, 7.669, 7.771, 7.805, 7.827, 7.867, 7.891, 7.925, 7.979, 7.999, 8.041, 8.081, 8.095, 8.135, 8.205, 8.253, 8.309, 8.425, 8.453, 8.473, 8.545, 8.581, 8.663, 8.697, 8.771, 8.969, 9.063, 9.111, 9.167, 9.197, 9.177, 9.151, 9.211, 9.287, 9.313, 9.345, 9.487, 9.627, 9.673, 9.685, 9.705, 9.793, 9.929, 10.069, 10.329, 10.365, 10.457, 10.425, 10.385, 10.221, 10.201, 10.181, 10.581, 11.009, 11.009, 11.061, 11.181, 11.333, 11.437, 11.506, 11.536, 11.556, 11.599, 11.606, 11.606, 6.102, 6.122, 6.149, 6.195, 6.272, 6.302, 6.35, 6.445, 6.517, 6.609, 6.721, 6.746, 6.758, 6.795, 6.881, 6.978, 7.036, 7.119, 7.187, 7.227, 7.283, 7.303, 7.331, 7.351, 7.415, 7.453, 7.469, 7.569, 7.685, 7.749, 7.825, 7.867, 7.917, 7.937, 7.915, 8.037, 8.045, 8.185, 8.289, 8.351, 8.442, 8.499, 8.529, 8.583, 8.667, 8.841, 8.97, 9.0, 9.024, 9.114, 9.228, 9.396, 9.537, 9.645, 9.693, 9.753, 9.807, 9.927, 10.272, 10.335, 10.44, 10.122, 10.356, 10.182, 10.206, 10.344, 10.986, 10.986, 11.124, 11.148, 11.412, 11.394}
    temp_qc = 
      {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
    cndc = 
      {3.72344, 3.86723, 3.9826, 4.13482, 4.22476, 3.65783, 3.66195, 3.66572, 3.66709, 3.66968, 3.67219, 3.67275, 3.67334, 3.67356, 3.6738, 3.67401, 3.67433, 3.67438, 3.67513, 3.67512, 3.67525, 3.6759, 3.67543, 3.67498, 3.67475, 3.67439, 3.67318, 3.67311, 3.67293, 3.67383, 3.67412, 3.67431, 3.67094, 3.65833, 3.64855, 3.65002, 3.64905, 3.65236, 3.6567, 3.65915, 3.66303, 3.66999, 3.67475, 3.67626, 3.67731, 3.6796, 3.68218, 3.6844, 3.68828, 3.69187, 3.693, 3.69486, 3.694, 3.69443, 3.6945, 3.69008, 3.69077, 3.68443, 3.66452, 3.64999, 3.64981, 3.63718, 3.66458, 3.68168, 3.68856, 3.68274, 3.67509, 3.67383, 3.67327, 3.67168, 3.6705, 3.66979, 3.66953, 3.66928, 3.66923, 3.66917, 3.66909, 3.66893, 3.66793, 3.66523, 3.66469, 3.66505, 3.66587, 3.66748, 3.67014, 3.67076, 3.67284, 3.67349, 3.674, 3.67429, 3.67526, 3.67651, 3.67759, 3.67975, 3.68021, 3.67988, 3.67987, 3.68101, 3.68509, 3.68521, 3.68415, 3.66857, 3.66883, 3.66907, 3.66939, 3.66972, 3.67006, 3.67011, 3.67061, 3.6713, 3.67261, 3.67423, 3.67551, 3.6756, 3.67536, 3.67538, 3.67675, 3.67879, 3.68126, 3.68248, 3.68106, 3.67104, 3.66548, 3.65582, 3.65614, 3.65275, 3.65229, 3.65254, 3.6513, 3.64995, 3.65023, 3.65057, 3.65143, 3.65154, 3.65209, 3.65376, 3.65754, 3.65829, 3.65903, 3.65993, 3.66544, 3.67239, 3.6798, 3.68705, 3.69045, 3.69386, 3.69477, 3.69034, 3.68221, 3.68158, 3.67665, 3.65765, 3.64265, 3.63962, 3.63433, 3.63226, 3.64036, 3.66498, 3.67592, 3.68383, 3.68374, 3.67901, 3.67437, 3.67274, 3.67146, 3.67067, 3.67002, 3.66992, 3.668, 3.66637, 3.66529, 3.6656, 3.66761, 3.66832, 3.66957, 3.67445, 3.67952, 3.68449, 3.68731, 3.68763, 3.68865, 3.68915, 3.6897, 3.6908, 3.6912, 3.69392, 3.69288, 3.69443, 3.69484, 3.6955, 3.66724, 3.66741, 3.66766, 3.6688, 3.67245, 3.67428, 3.67478, 3.67556, 3.67606, 3.67597, 3.67616, 3.67664, 3.67696, 3.67743, 3.67821, 3.6789, 3.67978, 3.68236, 3.68349, 3.68059, 3.67324, 3.66777, 3.65823, 3.65424, 3.65161, 3.65005, 3.64979, 3.64925, 3.64851, 3.64817, 3.64755, 3.64754, 3.64757, 3.64955, 3.65354, 3.65477, 3.6585, 3.66159, 3.67217, 3.68688, 3.68848, 3.6907, 3.6941, 3.69613, 3.6958, 3.69184, 3.67874, 3.66901, 3.65894, 3.65285, 3.65085, 3.64937, 3.64884, 3.64841, 3.64835, 3.64831, 3.64758, 3.63858, 3.6299, 3.63014, 3.62999, 3.63068, 3.65467, 3.6691, 3.67753, 3.67767, 3.67343, 3.6696, 3.66864, 3.66689, 3.66573, 3.66594, 3.66674, 3.66788, 3.67477, 3.68132, 3.68315, 3.68517, 3.68616, 3.68843, 3.68947, 3.69116, 3.69127, 3.69265, 3.69429, 3.69524, 3.69638, 3.69817, 3.69922, 3.67777, 3.67774, 3.67715, 3.6764, 3.67535, 3.67941, 3.68038, 3.6819, 3.68221, 3.67711, 3.67046, 3.66652, 3.66369, 3.66083, 3.65881, 3.65766, 3.65723, 3.65453, 3.65251, 3.65081, 3.65015, 3.65012, 3.65037, 3.65095, 3.65393, 3.65476, 3.65594, 3.6565, 3.65751, 3.65809, 3.66003, 3.66128, 3.66192, 3.66106, 3.66078, 3.66191, 3.66277, 3.66422, 3.67259, 3.68519, 3.69297, 3.69526, 3.69132, 3.68249, 3.67514, 3.67174, 3.66363, 3.65785, 3.6587, 3.65988, 3.66038, 3.66712, 3.66282, 3.65308, 3.65639, 3.69234, 3.6869, 3.68649, 3.68567, 3.68432, 3.68383, 3.68623, 3.68714, 3.68422, 3.68085, 3.67853, 3.6773, 3.67628, 3.67544, 3.6725, 3.67121, 3.67041, 3.66851, 3.66671, 3.66626, 3.66707, 3.67161, 3.67679, 3.682, 3.68573, 3.68626, 3.68605, 3.68682, 3.68713, 3.68842, 3.68883, 3.69098, 3.69155, 3.69438, 3.69681, 3.69739, 3.69888, 3.70367, 3.67307, 3.67305, 3.67315, 3.6734, 3.67229, 3.67184, 3.67151, 3.67043, 3.67039, 3.66912, 3.6686, 3.6667, 3.66665, 3.66568, 3.66469, 3.66164, 3.65984, 3.65826, 3.65689, 3.65614, 3.65588, 3.65555, 3.65518, 3.65512, 3.65505, 3.65479, 3.65422, 3.65433, 3.65427, 3.65456, 3.65642, 3.66338, 3.66902, 3.67092, 3.67237, 3.6748, 3.67755, 3.68354, 3.69506, 3.69543, 3.69551, 3.69442, 3.68754, 3.67731, 3.66621, 3.66687, 3.67977, 3.68216, 3.68602, 3.68778, 3.68984, 3.70015, 3.69758, 3.69176, 3.68963, 3.68789, 3.68715, 3.68438, 3.68206, 3.67773, 3.67608, 3.67583, 3.67477, 3.67533, 3.67418, 3.67342, 3.67215, 3.67015, 3.66957, 3.66844, 3.66756, 3.66805, 3.67147, 3.67598, 3.68113, 3.68354, 3.68572, 3.68833, 3.68928, 3.68949, 3.68972, 3.6903, 3.69098, 3.69267, 3.69578, 3.6969, 3.69817, 3.69921, 3.69987, 3.70549, 3.71379, 3.62466, 3.62489, 3.62493, 3.62487, 3.62499, 3.62464, 3.62464, 3.62428, 3.62418, 3.62422, 3.62426, 3.6353, 3.64716, 3.65186, 3.65209, 3.66081, 3.66465, 3.66532, 3.66761, 3.66903, 3.66926, 3.67039, 3.67169, 3.67224, 3.67096, 3.66547, 3.66056, 3.65879, 3.65655, 3.65621, 3.65567, 3.65559, 3.65687, 3.67613, 3.67974, 3.68077, 3.68651, 3.69257, 3.67872, 3.67127, 3.66644, 3.671, 3.69729, 3.69375, 3.67882, 3.67591, 3.67473, 3.66988, 3.6713, 3.67517, 3.68214, 3.68364, 3.6854, 3.688, 3.68882, 3.68959, 3.69339, 3.6978, 3.70464, 3.71426, 3.61275, 3.61279, 3.61292, 3.61276, 3.61307, 3.6129, 3.61318, 3.61264, 3.614, 3.61629, 3.61695, 3.61737, 3.61695, 3.61662, 3.6162, 3.61698, 3.62392, 3.62715, 3.64083, 3.65135, 3.65387, 3.65656, 3.65914, 3.66292, 3.66586, 3.6673, 3.67144, 3.66944, 3.66481, 3.66313, 3.65793, 3.65749, 3.65695, 3.6565, 3.65693, 3.66955, 3.68305, 3.68793, 3.68844, 3.68866, 3.69002, 3.69101, 3.6871, 3.6806, 3.67729, 3.6585, 3.67454, 3.68338, 3.67454, 3.67469, 3.67845, 3.68814, 3.69099, 3.69142, 3.69023, 3.68952, 3.68893, 3.68977, 3.69014, 3.69112, 3.69713, 3.69918, 3.70377, 3.71652, 3.60583, 3.60596, 3.60599, 3.60619, 3.6063, 3.60695, 3.60687, 3.60805, 3.60993, 3.61214, 3.61431, 3.61773, 3.62616, 3.63438, 3.63755, 3.64162, 3.64669, 3.65047, 3.65677, 3.65992, 3.66045, 3.66144, 3.66744, 3.6699, 3.67019, 3.6698, 3.66869, 3.66695, 3.66507, 3.66214, 3.66029, 3.65864, 3.65775, 3.65723, 3.65966, 3.66637, 3.6735, 3.67867, 3.68169, 3.6845, 3.68564, 3.68522, 3.68281, 3.65936, 3.65133, 3.66522, 3.6726, 3.66985, 3.67161, 3.67417, 3.67855, 3.69163, 3.6969, 3.69773, 3.69804, 3.69807, 3.69789, 3.6982, 3.69878, 3.70267, 3.71489, 3.71593, 3.56861, 3.57101, 3.57194, 3.5727, 3.57363, 3.57545, 3.57655, 3.57691, 3.57835, 3.57976, 3.58091, 3.58208, 3.58351, 3.5863, 3.58791, 3.58952, 3.59349, 3.59546, 3.59716, 3.60013, 3.60344, 3.60839, 3.61387, 3.61638, 3.6199, 3.6345, 3.64083, 3.64538, 3.64755, 3.64963, 3.65188, 3.65377, 3.65837, 3.66043, 3.66149, 3.66239, 3.66456, 3.6667, 3.66717, 3.66542, 3.66417, 3.66307, 3.66143, 3.66075, 3.65987, 3.65918, 3.65848, 3.65952, 3.66563, 3.67619, 3.6784, 3.68144, 3.68318, 3.68335, 3.68084, 3.6683, 3.63942, 3.63792, 3.64935, 3.66925, 3.66352, 3.66864, 3.67407, 3.68427, 3.70219, 3.70506, 3.70645, 3.70818, 3.7097, 3.71061, 3.71032, 3.71095, 3.712, 3.71824, 3.72213, 3.72292, 3.72311, 3.53943, 3.53974, 3.54096, 3.54171, 3.54191, 3.54202, 3.54194, 3.54312, 3.54701, 3.55604, 3.56289, 3.56795, 3.57138, 3.57389, 3.57677, 3.57955, 3.58061, 3.58084, 3.58199, 3.58405, 3.59081, 3.59377, 3.59419, 3.5964, 3.59789, 3.59932, 3.6019, 3.60394, 3.60598, 3.6092, 3.61126, 3.62194, 3.63374, 3.63909, 3.64426, 3.64854, 3.65451, 3.65792, 3.65988, 3.66166, 3.66404, 3.66507, 3.66548, 3.66581, 3.66664, 3.66968, 3.66972, 3.66901, 3.6685, 3.66696, 3.66663, 3.66452, 3.66277, 3.65484, 3.65064, 3.65196, 3.66502, 3.67488, 3.68169, 3.68367, 3.67825, 3.66471, 3.65542, 3.65253, 3.64, 3.65739, 3.67333, 3.67732, 3.67758, 3.68014, 3.68384, 3.69749, 3.70636, 3.71308, 3.71731, 3.72338, 3.7272, 3.72783, 3.72854, 3.72977, 3.73207, 3.73271, 3.73297, 3.73319, 3.54902, 3.54996, 3.55344, 3.55627, 3.55702, 3.55793, 3.55993, 3.56336, 3.56733, 3.57138, 3.57317, 3.57507, 3.57552, 3.57659, 3.57757, 3.57965, 3.58534, 3.59157, 3.59708, 3.60097, 3.60557, 3.60827, 3.61033, 3.61112, 3.61081, 3.61042, 3.61067, 3.61145, 3.61195, 3.62609, 3.63298, 3.63878, 3.6424, 3.64365, 3.64452, 3.64813, 3.65561, 3.65667, 3.65851, 3.65975, 3.66179, 3.66461, 3.66727, 3.66929, 3.67195, 3.67242, 3.67353, 3.67429, 3.67243, 3.66199, 3.64068, 3.63545, 3.63734, 3.64952, 3.65897, 3.66409, 3.67726, 3.68535, 3.68634, 3.68291, 3.67812, 3.67071, 3.65374, 3.64722, 3.63875, 3.63709, 3.64282, 3.64954, 3.68462, 3.68502, 3.68231, 3.68228, 3.69738, 3.71241, 3.71633, 3.71747, 3.71748, 3.71626, 3.71467, 3.71272, 3.71121, 3.71908, 3.72125, 3.72065, 3.56175, 3.56678, 3.5709, 3.57228, 3.57621, 3.57885, 3.57921, 3.5793, 3.58091, 3.58396, 3.58522, 3.58875, 3.59055, 3.59163, 3.59505, 3.59875, 3.60408, 3.60816, 3.6095, 3.61003, 3.61319, 3.61272, 3.61516, 3.61884, 3.626, 3.62844, 3.62879, 3.62931, 3.63038, 3.6319, 3.63242, 3.63827, 3.64125, 3.64366, 3.64517, 3.64605, 3.64721, 3.64963, 3.65531, 3.65745, 3.6586, 3.65931, 3.66001, 3.66213, 3.66478, 3.66557, 3.66977, 3.67232, 3.67319, 3.67414, 3.67482, 3.67534, 3.67586, 3.67578, 3.64579, 3.63521, 3.63518, 3.64165, 3.65322, 3.67827, 3.68687, 3.68395, 3.67562, 3.64567, 3.62834, 3.62839, 3.63919, 3.64674, 3.65139, 3.66979, 3.67221, 3.69416, 3.68496, 3.68706, 3.69205, 3.69751, 3.70552, 3.71062, 3.7128, 3.71311, 3.71301, 3.71491, 3.71802, 3.71916, 3.71961, 3.71979, 3.71927, 3.49824, 3.5042, 3.51094, 3.51259, 3.51517, 3.51826, 3.52344, 3.52672, 3.53045, 3.53627, 3.53784, 3.54112, 3.54368, 3.54615, 3.5486, 3.54971, 3.55922, 3.56623, 3.56943, 3.57753, 3.58118, 3.58991, 3.59684, 3.60068, 3.60679, 3.62294, 3.63264, 3.63679, 3.64027, 3.64249, 3.64557, 3.6485, 3.65476, 3.65775, 3.66364, 3.6683, 3.67286, 3.67553, 3.67763, 3.67835, 3.64454, 3.65232, 3.66067, 3.65032, 3.6283, 3.65736, 3.67821, 3.66128, 3.69021, 3.69621, 3.69814, 3.70911, 3.71083, 3.7096, 3.71347, 3.71598, 3.71686, 3.71693, 3.48784, 3.4907, 3.49498, 3.49842, 3.50109, 3.50391, 3.50773, 3.50865, 3.50829, 3.50872, 3.51078, 3.5143, 3.52635, 3.53995, 3.54596, 3.54716, 3.5538, 3.55737, 3.56418, 3.56675, 3.57085, 3.57386, 3.57697, 3.57899, 3.58128, 3.58712, 3.59496, 3.60125, 3.61193, 3.62672, 3.63375, 3.63742, 3.64163, 3.64608, 3.65055, 3.6534, 3.6592, 3.66806, 3.67616, 3.68055, 3.68205, 3.677, 3.65837, 3.65732, 3.65732, 3.64252, 3.62551, 3.64748, 3.67402, 3.67058, 3.67119, 3.68853, 3.69122, 3.69493, 3.70898, 3.71436, 3.71598, 3.71404, 3.7126, 3.71195, 3.47926, 3.48301, 3.48315, 3.48813, 3.49289, 3.4932, 3.4938, 3.49593, 3.49696, 3.49944, 3.50174, 3.50809, 3.51003, 3.51378, 3.52077, 3.52678, 3.53505, 3.5476, 3.55645, 3.55813, 3.56244, 3.56837, 3.57212, 3.57334, 3.57548, 3.57661, 3.58099, 3.58458, 3.58618, 3.58884, 3.60068, 3.60765, 3.61853, 3.62915, 3.63465, 3.63779, 3.63823, 3.63987, 3.64608, 3.64912, 3.6591, 3.66789, 3.66985, 3.67371, 3.67672, 3.68355, 3.68641, 3.68831, 3.69067, 3.68373, 3.67125, 3.66253, 3.65898, 3.66606, 3.67395, 3.68035, 3.6921, 3.68432, 3.69007, 3.68715, 3.69643, 3.70249, 3.7036, 3.70494, 3.71, 3.71577, 3.7162, 3.71566, 3.71509, 3.46818, 3.46826, 3.46723, 3.46779, 3.47255, 3.47638, 3.47889, 3.48355, 3.48776, 3.49161, 3.49547, 3.4959, 3.49569, 3.49567, 3.49581, 3.49676, 3.49806, 3.49955, 3.50203, 3.5112, 3.51458, 3.51615, 3.52018, 3.52538, 3.53032, 3.53372, 3.5411, 3.54352, 3.54539, 3.54843, 3.55003, 3.55428, 3.5609, 3.56478, 3.56738, 3.57236, 3.5745, 3.5745, 3.58155, 3.58732, 3.59082, 3.60094, 3.6142, 3.62978, 3.63448, 3.63632, 3.63975, 3.64347, 3.64588, 3.65807, 3.66192, 3.66294, 3.66378, 3.6664, 3.67713, 3.69126, 3.69396, 3.69514, 3.68533, 3.66643, 3.66278, 3.66672, 3.66791, 3.67171, 3.67977, 3.68396, 3.66535, 3.6489, 3.67815, 3.69649, 3.69332, 3.70241, 3.70473, 3.70381, 3.70477, 3.70596, 3.70709, 3.70879, 3.71492, 3.71545, 3.44755, 3.44744, 3.4474, 3.44698, 3.44633, 3.44684, 3.44853, 3.45335, 3.45879, 3.46028, 3.46258, 3.46624, 3.47243, 3.47511, 3.47842, 3.48026, 3.4812, 3.48386, 3.48688, 3.48883, 3.49168, 3.49888, 3.51134, 3.51602, 3.52222, 3.52762, 3.53112, 3.53424, 3.538, 3.54167, 3.54244, 3.54458, 3.54834, 3.55331, 3.55808, 3.55942, 3.55995, 3.56091, 3.56242, 3.56793, 3.57208, 3.57222, 3.57462, 3.57713, 3.58254, 3.58906, 3.59367, 3.60162, 3.61328, 3.62359, 3.63625, 3.63871, 3.64072, 3.64178, 3.64254, 3.64582, 3.64875, 3.64973, 3.65936, 3.66784, 3.67416, 3.67694, 3.69033, 3.70228, 3.70683, 3.70819, 3.71191, 3.71549, 3.71385, 3.7061, 3.69909, 3.69294, 3.68281, 3.67164, 3.64512, 3.58477, 3.58548, 3.62294, 3.6423, 3.66992, 3.68271, 3.69458, 3.69574, 3.70134, 3.70486, 3.70499, 3.45254, 3.45359, 3.45731, 3.46075, 3.46098, 3.46219, 3.46442, 3.46845, 3.4713, 3.47263, 3.4745, 3.47493, 3.47635, 3.47867, 3.48081, 3.4843, 3.4868, 3.48903, 3.49099, 3.49269, 3.49745, 3.49995, 3.50463, 3.52036, 3.52894, 3.53162, 3.53322, 3.53625, 3.53811, 3.5406, 3.54472, 3.54612, 3.54915, 3.55162, 3.55174, 3.55431, 3.55998, 3.56337, 3.56805, 3.57877, 3.58138, 3.58298, 3.58856, 3.59114, 3.59736, 3.5992, 3.6047, 3.62258, 3.6304, 3.63382, 3.63788, 3.63888, 3.63386, 3.62955, 3.63251, 3.63753, 3.63979, 3.64262, 3.65407, 3.66388, 3.6668, 3.66749, 3.66852, 3.67167, 3.67901, 3.68867, 3.71033, 3.71403, 3.7195, 3.70525, 3.69782, 3.67159, 3.66405, 3.65413, 3.68168, 3.70787, 3.69437, 3.68655, 3.69211, 3.69931, 3.70472, 3.70839, 3.70886, 3.71038, 3.71428, 3.71499, 3.71482, 3.39513, 3.39674, 3.39858, 3.40203, 3.40809, 3.41036, 3.41405, 3.42152, 3.42729, 3.4345, 3.44388, 3.44588, 3.44669, 3.44967, 3.45653, 3.46447, 3.46935, 3.47632, 3.48175, 3.48511, 3.48973, 3.4912, 3.49311, 3.49404, 3.49877, 3.5019, 3.50303, 3.51196, 3.52225, 3.52699, 3.5332, 3.53492, 3.53821, 3.53896, 3.53468, 3.54515, 3.54518, 3.55664, 3.56531, 3.57027, 3.57825, 3.58304, 3.58499, 3.58856, 3.59515, 3.60996, 3.62134, 3.6212, 3.61973, 3.62621, 3.63449, 3.6485, 3.658, 3.66475, 3.66737, 3.67127, 3.67482, 3.68324, 3.70837, 3.70631, 3.71105, 3.66469, 3.66884, 3.63063, 3.62083, 3.62521, 3.68269, 3.66949, 3.6695, 3.66857, 3.69283, 3.69122}
    cndc_qc = 
      {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
    chla = 
      {0.228, 0.228, 0.231, 0.219, 0.216, 0.192, 0.189, 0.189, 0.195, 0.192, 0.192, 0.192, 0.189, 0.192, 0.189, 0.189, 0.192, 0.192, 0.195, 0.192, 0.192, 0.192, 0.189, 0.195, 0.192, 0.192, 0.198, 0.198, 0.195, 0.195, 0.192, 0.195, 0.198, 0.192, 0.198, 0.201, 0.198, 0.195, 0.198, 0.198, 0.201, 0.198, 0.201, 0.201, 0.201, 0.201, 0.198, 0.204, 0.198, 0.201, 0.198, 0.207, 0.207, 0.21, 0.216, 0.219, 0.222, 0.234, 0.243, 0.249, 0.288, 0.339, 0.366, 0.387, 0.408, 0.417, 0.408, 0.432, 0.435, 0.429, 0.42, 0.417, 0.405, 0.417, 0.426, 0.411, 0.438, 0.414, 0.42, 0.426, 0.429, 0.435, 0.426, 0.447, 0.435, 0.429, 0.45, 0.42, 0.432, 0.435, 0.426, 0.417, 0.396, 0.372, 0.351, 0.339, 0.318, 0.294, 0.285, 0.276, 0.276, 0.189, 0.186, 0.192, 0.189, 0.189, 0.195, 0.186, 0.192, 0.189, 0.189, 0.189, 0.189, 0.192, 0.192, 0.192, 0.192, 0.192, 0.195, 0.195, 0.192, 0.201, 0.195, 0.195, 0.195, 0.198, 0.195, 0.192, 0.195, 0.198, 0.195, 0.195, 0.195, 0.195, 0.201, 0.198, 0.198, 0.201, 0.198, 0.201, 0.198, 0.195, 0.195, 0.198, 0.195, 0.201, 0.201, 0.213, 0.21, 0.204, 0.216, 0.222, 0.234, 0.249, 0.261, 0.291, 0.33, 0.351, 0.375, 0.396, 0.396, 0.417, 0.402, 0.411, 0.408, 0.387, 0.384, 0.39, 0.39, 0.411, 0.417, 0.435, 0.456, 0.453, 0.456, 0.423, 0.411, 0.393, 0.366, 0.375, 0.36, 0.357, 0.345, 0.339, 0.312, 0.312, 0.291, 0.288, 0.276, 0.267, 0.192, 0.192, 0.186, 0.189, 0.189, 0.186, 0.192, 0.192, 0.189, 0.189, 0.189, 0.192, 0.192, 0.192, 0.189, 0.192, 0.192, 0.192, 0.189, 0.189, 0.189, 0.192, 0.195, 0.192, 0.192, 0.192, 0.192, 0.192, 0.189, 0.192, 0.195, 0.192, 0.195, 0.192, 0.192, 0.198, 0.198, 0.198, 0.195, 0.198, 0.198, 0.198, 0.201, 0.204, 0.198, 0.204, 0.21, 0.213, 0.222, 0.216, 0.222, 0.225, 0.222, 0.216, 0.219, 0.222, 0.228, 0.246, 0.273, 0.273, 0.27, 0.294, 0.333, 0.354, 0.369, 0.378, 0.411, 0.375, 0.402, 0.39, 0.408, 0.423, 0.462, 0.462, 0.444, 0.423, 0.414, 0.378, 0.375, 0.366, 0.351, 0.324, 0.315, 0.297, 0.288, 0.276, 0.27, 0.255, 0.258, 0.192, 0.186, 0.192, 0.189, 0.186, 0.192, 0.189, 0.189, 0.189, 0.195, 0.192, 0.192, 0.186, 0.189, 0.186, 0.192, 0.192, 0.189, 0.195, 0.192, 0.192, 0.189, 0.192, 0.192, 0.189, 0.192, 0.192, 0.192, 0.189, 0.189, 0.192, 0.195, 0.192, 0.192, 0.195, 0.195, 0.195, 0.192, 0.192, 0.195, 0.192, 0.198, 0.198, 0.201, 0.204, 0.207, 0.213, 0.219, 0.237, 0.231, 0.231, 0.243, 0.249, 0.255, 0.318, 0.333, 0.327, 0.339, 0.339, 0.351, 0.381, 0.39, 0.381, 0.39, 0.381, 0.399, 0.381, 0.396, 0.426, 0.39, 0.396, 0.405, 0.408, 0.426, 0.447, 0.48, 0.474, 0.438, 0.42, 0.411, 0.429, 0.405, 0.387, 0.384, 0.363, 0.327, 0.312, 0.294, 0.288, 0.273, 0.273, 0.261, 0.252, 0.189, 0.186, 0.186, 0.189, 0.186, 0.186, 0.186, 0.192, 0.189, 0.189, 0.189, 0.186, 0.189, 0.192, 0.189, 0.189, 0.192, 0.192, 0.189, 0.192, 0.192, 0.192, 0.195, 0.189, 0.192, 0.192, 0.189, 0.192, 0.192, 0.192, 0.192, 0.192, 0.192, 0.195, 0.195, 0.198, 0.195, 0.195, 0.195, 0.195, 0.198, 0.201, 0.204, 0.213, 0.222, 0.231, 0.264, 0.276, 0.279, 0.279, 0.318, 0.354, 0.366, 0.378, 0.39, 0.384, 0.396, 0.402, 0.405, 0.429, 0.42, 0.405, 0.432, 0.414, 0.417, 0.402, 0.411, 0.417, 0.423, 0.459, 0.474, 0.474, 0.438, 0.45, 0.426, 0.417, 0.417, 0.426, 0.417, 0.396, 0.396, 0.381, 0.369, 0.318, 0.309, 0.3, 0.288, 0.276, 0.267, 0.252, 0.249, 0.192, 0.192, 0.192, 0.192, 0.189, 0.189, 0.192, 0.192, 0.192, 0.192, 0.192, 0.189, 0.192, 0.189, 0.189, 0.192, 0.189, 0.189, 0.192, 0.192, 0.189, 0.189, 0.189, 0.189, 0.189, 0.192, 0.189, 0.189, 0.192, 0.192, 0.192, 0.189, 0.189, 0.195, 0.195, 0.192, 0.195, 0.198, 0.207, 0.21, 0.213, 0.237, 0.318, 0.363, 0.408, 0.426, 0.42, 0.45, 0.447, 0.441, 0.405, 0.408, 0.42, 0.417, 0.429, 0.405, 0.357, 0.312, 0.288, 0.264, 0.192, 0.192, 0.189, 0.192, 0.189, 0.192, 0.192, 0.192, 0.189, 0.192, 0.189, 0.189, 0.192, 0.192, 0.189, 0.192, 0.192, 0.189, 0.189, 0.189, 0.189, 0.186, 0.192, 0.189, 0.186, 0.189, 0.192, 0.189, 0.192, 0.189, 0.189, 0.192, 0.189, 0.189, 0.189, 0.192, 0.195, 0.195, 0.198, 0.195, 0.198, 0.198, 0.201, 0.204, 0.207, 0.225, 0.294, 0.354, 0.378, 0.378, 0.393, 0.39, 0.396, 0.399, 0.396, 0.399, 0.405, 0.414, 0.426, 0.423, 0.396, 0.348, 0.309, 0.291, 0.189, 0.192, 0.189, 0.189, 0.192, 0.189, 0.192, 0.192, 0.192, 0.189, 0.189, 0.192, 0.189, 0.189, 0.189, 0.189, 0.192, 0.189, 0.189, 0.189, 0.192, 0.189, 0.189, 0.186, 0.189, 0.189, 0.186, 0.192, 0.189, 0.189, 0.189, 0.189, 0.189, 0.192, 0.189, 0.192, 0.192, 0.192, 0.192, 0.195, 0.195, 0.198, 0.198, 0.219, 0.273, 0.306, 0.336, 0.351, 0.366, 0.372, 0.414, 0.396, 0.405, 0.399, 0.399, 0.399, 0.393, 0.39, 0.39, 0.375, 0.354, 0.33, 0.192, 0.189, 0.192, 0.192, 0.189, 0.192, 0.192, 0.192, 0.195, 0.192, 0.192, 0.192, 0.192, 0.192, 0.192, 0.192, 0.192, 0.195, 0.189, 0.189, 0.189, 0.192, 0.192, 0.189, 0.189, 0.192, 0.192, 0.192, 0.192, 0.189, 0.189, 0.096, 0.189, 0.189, 0.189, 0.186, 0.192, 0.189, 0.192, 0.189, 0.189, 0.192, 0.189, 0.186, 0.189, 0.189, 0.189, 0.192, 0.192, 0.192, 0.195, 0.195, 0.195, 0.198, 0.198, 0.207, 0.237, 0.249, 0.288, 0.318, 0.339, 0.375, 0.408, 0.423, 0.456, 0.447, 0.45, 0.447, 0.435, 0.435, 0.42, 0.405, 0.396, 0.381, 0.369, 0.363, 0.363, 0.195, 0.195, 0.195, 0.195, 0.195, 0.195, 0.195, 0.195, 0.195, 0.195, 0.195, 0.192, 0.195, 0.198, 0.192, 0.195, 0.195, 0.195, 0.192, 0.195, 0.195, 0.195, 0.192, 0.195, 0.195, 0.195, 0.195, 0.195, 0.195, 0.192, 0.192, 0.192, 0.192, 0.192, 0.192, 0.192, 0.192, 0.192, 0.186, 0.192, 0.192, 0.189, 0.189, 0.189, 0.189, 0.192, 0.189, 0.192, 0.192, 0.192, 0.189, 0.192, 0.189, 0.189, 0.195, 0.192, 0.195, 0.192, 0.195, 0.195, 0.198, 0.201, 0.21, 0.213, 0.231, 0.291, 0.378, 0.399, 0.408, 0.414, 0.423, 0.414, 0.417, 0.423, 0.411, 0.411, 0.408, 0.372, 0.348, 0.372, 0.375, 0.378, 0.378, 0.378, 0.192, 0.192, 0.192, 0.195, 0.192, 0.192, 0.195, 0.192, 0.192, 0.192, 0.192, 0.192, 0.195, 0.192, 0.192, 0.195, 0.192, 0.195, 0.192, 0.192, 0.189, 0.192, 0.192, 0.192, 0.192, 0.189, 0.189, 0.192, 0.192, 0.192, 0.189, 0.189, 0.192, 0.189, 0.192, 0.192, 0.189, 0.189, 0.189, 0.189, 0.189, 0.189, 0.189, 0.189, 0.189, 0.192, 0.189, 0.189, 0.186, 0.189, 0.192, 0.192, 0.192, 0.189, 0.198, 0.192, 0.195, 0.195, 0.198, 0.198, 0.195, 0.201, 0.201, 0.21, 0.219, 0.231, 0.255, 0.297, 0.396, 0.423, 0.432, 0.417, 0.393, 0.363, 0.366, 0.369, 0.36, 0.357, 0.345, 0.348, 0.333, 0.297, 0.294, 0.297, 0.192, 0.192, 0.189, 0.186, 0.189, 0.189, 0.189, 0.189, 0.192, 0.189, 0.192, 0.189, 0.189, 0.189, 0.189, 0.192, 0.189, 0.189, 0.192, 0.189, 0.186, 0.189, 0.189, 0.189, 0.189, 0.189, 0.189, 0.186, 0.192, 0.189, 0.189, 0.189, 0.189, 0.186, 0.189, 0.189, 0.189, 0.192, 0.189, 0.189, 0.189, 0.189, 0.186, 0.189, 0.189, 0.186, 0.189, 0.189, 0.189, 0.189, 0.186, 0.189, 0.189, 0.189, 0.189, 0.192, 0.189, 0.192, 0.189, 0.192, 0.198, 0.192, 0.195, 0.21, 0.219, 0.231, 0.246, 0.255, 0.273, 0.288, 0.276, 0.312, 0.336, 0.336, 0.369, 0.372, 0.369, 0.36, 0.348, 0.321, 0.309, 0.3, 0.288, 0.3, 0.288, 0.288, 0.285, 0.195, 0.195, 0.198, 0.195, 0.198, 0.198, 0.198, 0.198, 0.195, 0.198, 0.195, 0.198, 0.198, 0.198, 0.195, 0.195, 0.195, 0.195, 0.192, 0.195, 0.195, 0.192, 0.195, 0.192, 0.192, 0.192, 0.192, 0.192, 0.189, 0.192, 0.192, 0.189, 0.189, 0.189, 0.189, 0.189, 0.189, 0.189, 0.189, 0.186, 0.189, 0.189, 0.192, 0.198, 0.225, 0.264, 0.267, 0.261, 0.189, 0.318, 0.357, 0.333, 0.324, 0.327, 0.288, 0.285, 0.279, 0.279, 0.195, 0.195, 0.198, 0.195, 0.195, 0.195, 0.198, 0.195, 0.198, 0.195, 0.195, 0.195, 0.195, 0.195, 0.198, 0.195, 0.195, 0.198, 0.195, 0.192, 0.192, 0.192, 0.192, 0.192, 0.192, 0.192, 0.189, 0.192, 0.192, 0.189, 0.189, 0.189, 0.189, 0.189, 0.192, 0.192, 0.192, 0.189, 0.189, 0.192, 0.192, 0.189, 0.189, 0.192, 0.192, 0.195, 0.198, 0.264, 0.279, 0.267, 0.267, 0.297, 0.33, 0.366, 0.33, 0.315, 0.318, 0.3, 0.3, 0.303, 0.198, 0.198, 0.198, 0.198, 0.198, 0.198, 0.198, 0.198, 0.198, 0.198, 0.198, 0.198, 0.198, 0.198, 0.198, 0.195, 0.195, 0.195, 0.198, 0.195, 0.195, 0.195, 0.195, 0.195, 0.192, 0.195, 0.192, 0.192, 0.192, 0.195, 0.192, 0.192, 0.192, 0.192, 0.189, 0.192, 0.192, 0.192, 0.192, 0.189, 0.192, 0.189, 0.189, 0.189, 0.189, 0.189, 0.192, 0.201, 0.189, 0.192, 0.195, 0.195, 0.198, 0.204, 0.213, 0.222, 0.243, 0.291, 0.297, 0.351, 0.339, 0.321, 0.321, 0.318, 0.318, 0.297, 0.297, 0.288, 0.291, 0.201, 0.201, 0.198, 0.204, 0.201, 0.198, 0.201, 0.201, 0.198, 0.201, 0.198, 0.201, 0.201, 0.201, 0.201, 0.198, 0.201, 0.201, 0.201, 0.198, 0.198, 0.198, 0.198, 0.195, 0.198, 0.198, 0.198, 0.195, 0.198, 0.198, 0.195, 0.195, 0.198, 0.195, 0.195, 0.198, 0.195, 0.195, 0.192, 0.195, 0.195, 0.192, 0.195, 0.195, 0.192, 0.192, 0.192, 0.189, 0.192, 0.192, 0.192, 0.189, 0.189, 0.189, 0.192, 0.192, 0.189, 0.192, 0.195, 0.195, 0.198, 0.198, 0.204, 0.21, 0.21, 0.216, 0.222, 0.228, 0.255, 0.291, 0.333, 0.318, 0.327, 0.333, 0.33, 0.33, 0.324, 0.318, 0.315, 0.312, 0.201, 0.201, 0.201, 0.201, 0.201, 0.201, 0.201, 0.198, 0.201, 0.201, 0.198, 0.201, 0.198, 0.198, 0.198, 0.201, 0.198, 0.201, 0.198, 0.198, 0.198, 0.198, 0.198, 0.198, 0.198, 0.195, 0.195, 0.195, 0.195, 0.195, 0.195, 0.195, 0.195, 0.195, 0.195, 0.195, 0.198, 0.195, 0.192, 0.195, 0.195, 0.192, 0.192, 0.195, 0.192, 0.195, 0.195, 0.192, 0.189, 0.189, 0.192, 0.192, 0.189, 0.195, 0.192, 0.192, 0.192, 0.192, 0.192, 0.192, 0.192, 0.192, 0.192, 0.192, 0.189, 0.192, 0.192, 0.192, 0.192, 0.195, 0.195, 0.198, 0.195, 0.198, 0.21, 0.216, 0.222, 0.249, 0.27, 0.306, 0.342, 0.366, 0.363, 0.339, 0.324, 0.321, 0.201, 0.198, 0.201, 0.201, 0.198, 0.198, 0.201, 0.198, 0.201, 0.198, 0.198, 0.198, 0.201, 0.198, 0.198, 0.198, 0.195, 0.198, 0.198, 0.195, 0.198, 0.198, 0.198, 0.198, 0.198, 0.195, 0.195, 0.195, 0.195, 0.195, 0.195, 0.195, 0.195, 0.195, 0.195, 0.195, 0.195, 0.195, 0.195, 0.195, 0.195, 0.195, 0.192, 0.195, 0.192, 0.192, 0.192, 0.192, 0.192, 0.192, 0.192, 0.192, 0.192, 0.189, 0.189, 0.189, 0.189, 0.189, 0.189, 0.192, 0.186, 0.189, 0.189, 0.189, 0.189, 0.189, 0.192, 0.195, 0.192, 0.192, 0.195, 0.195, 0.198, 0.201, 0.21, 0.231, 0.267, 0.312, 0.327, 0.321, 0.312, 0.309, 0.3, 0.294, 0.279, 0.27, 0.276, 0.201, 0.204, 0.201, 0.201, 0.201, 0.201, 0.201, 0.201, 0.201, 0.201, 0.201, 0.201, 0.201, 0.198, 0.201, 0.201, 0.198, 0.198, 0.201, 0.198, 0.198, 0.198, 0.198, 0.195, 0.198, 0.195, 0.195, 0.198, 0.195, 0.195, 0.195, 0.195, 0.192, 0.198, 0.195, 0.195, 0.195, 0.192, 0.192, 0.192, 0.192, 0.192, 0.192, 0.192, 0.192, 0.189, 0.189, 0.189, 0.189, 0.189, 0.189, 0.189, 0.189, 0.189, 0.189, 0.189, 0.189, 0.189, 0.189, 0.192, 0.192, 0.195, 0.195, 0.201, 0.213, 0.231, 0.285, 0.321, 0.339, 0.366, 0.342, 0.345}
    chla_qc = 
      {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
    doxy = 
      {281.3286, 271.566, 266.1686, 259.3934, 253.1995, 150.1627, 140.7665, 135.0039, 130.2885, 127.3307, 125.591, 124.3805, 123.7724, 123.3152, 123.0861, 122.9296, 122.929, 123.0763, 123.4629, 123.8468, 124.6823, 125.5296, 126.9756, 128.3544, 129.6549, 130.795, 131.9358, 133.0729, 134.2894, 135.2011, 135.9598, 137.0258, 139.2367, 143.3063, 149.2002, 153.3528, 156.6391, 160.4197, 162.6497, 164.262, 166.7454, 168.2479, 169.4996, 170.7171, 171.8571, 172.3524, 172.6611, 172.8945, 173.3745, 174.0123, 175.1756, 177.6312, 179.3946, 181.0844, 184.5439, 187.4522, 190.5378, 194.613, 200.6862, 205.0068, 211.314, 218.0895, 225.0267, 232.0703, 240.4886, 249.6433, 254.9023, 258.5113, 262.6507, 264.4027, 265.6957, 267.22, 267.7415, 268.1884, 268.5602, 268.9269, 269.0725, 269.2179, 269.5138, 269.6899, 269.9382, 270.261, 270.6453, 270.9841, 271.4468, 271.7552, 272.2398, 272.3525, 272.5074, 272.6175, 272.9359, 272.8293, 272.7203, 272.9521, 272.9895, 273.0543, 273.0366, 272.5531, 272.64, 272.7693, 272.5479, 123.8221, 122.3376, 121.3076, 120.7356, 120.3916, 120.0837, 119.9687, 119.8513, 119.8517, 120.2371, 120.9364, 121.8966, 123.9013, 125.5491, 127.1879, 128.4889, 130.1311, 130.9716, 132.112, 133.7878, 136.6202, 140.0444, 143.0572, 145.6763, 148.0845, 150.4063, 152.2343, 153.8013, 156.2503, 157.8634, 159.5815, 160.8051, 161.6016, 162.7053, 163.7096, 164.7795, 165.8459, 166.4472, 166.9844, 168.3318, 169.3402, 170.0664, 171.2495, 172.0933, 173.2803, 175.4242, 178.5603, 181.8317, 185.5739, 189.9827, 194.6092, 200.562, 206.3492, 212.0908, 216.6283, 222.0206, 227.4092, 231.8155, 239.1746, 245.5246, 251.0385, 256.5952, 260.1976, 262.4871, 264.7747, 265.9868, 266.9025, 267.6644, 268.2062, 268.5243, 269.2481, 270.0543, 270.4398, 271.0056, 271.0267, 271.0656, 271.0107, 271.208, 271.1895, 271.3369, 271.6351, 271.6213, 271.8897, 271.8362, 272.1856, 272.2055, 272.2859, 272.307, 272.378, 122.5643, 121.2323, 120.2047, 119.7924, 120.159, 120.8198, 121.5447, 122.6661, 124.2454, 125.9661, 127.3039, 128.5998, 129.6647, 130.5817, 131.2643, 131.7179, 132.0557, 132.2037, 132.9246, 134.1007, 135.8881, 138.705, 141.6878, 144.8117, 148.8915, 151.1456, 152.6275, 154.3765, 155.6284, 156.3817, 157.33, 158.1277, 159.0542, 160.9176, 162.3231, 163.4398, 165.3792, 166.3908, 167.9314, 169.4915, 170.2451, 171.1617, 172.0176, 173.7314, 175.6612, 178.3756, 183.4135, 187.6454, 191.5726, 195.8681, 198.8553, 200.7639, 202.7442, 203.7994, 204.3995, 205.0752, 206.2106, 209.5646, 214.8305, 219.1166, 221.9368, 224.2956, 228.8346, 233.9008, 242.4692, 248.9811, 254.5714, 258.4826, 261.933, 263.9141, 265.761, 267.1654, 268.1092, 269.0617, 269.5303, 269.7636, 270.0544, 270.856, 270.7017, 271.0114, 271.1573, 271.5409, 271.7172, 271.8687, 271.8679, 272.1658, 272.2362, 272.2021, 272.4237, 129.299, 128.4255, 128.4401, 129.4024, 130.3286, 131.3343, 132.0574, 132.5546, 133.6214, 135.2632, 137.583, 139.4832, 141.1173, 142.7946, 144.2033, 145.6836, 147.3537, 148.5327, 150.2456, 151.5445, 152.8066, 154.152, 155.265, 156.1382, 157.0351, 157.8749, 158.6799, 159.2871, 159.7461, 160.4277, 161.0164, 161.7119, 162.8207, 163.5382, 164.4517, 165.1842, 165.8815, 166.9945, 167.5557, 168.4155, 169.5262, 171.4859, 173.985, 179.0963, 182.8537, 185.7645, 190.1473, 193.3003, 196.767, 199.6111, 201.53, 205.5599, 208.8691, 211.4767, 215.7616, 222.2434, 226.2151, 230.4112, 233.962, 236.575, 240.1998, 244.9499, 248.3363, 251.8326, 256.1145, 258.8111, 260.9589, 262.5682, 264.4087, 265.5687, 266.369, 267.2067, 267.902, 268.2957, 269.0253, 269.5083, 270.2003, 270.0693, 270.5632, 271.0107, 271.1275, 271.3217, 271.8146, 271.8385, 272.0671, 272.2902, 272.3127, 272.3466, 272.4284, 272.6286, 272.7363, 272.6578, 272.4112, 136.5919, 135.4483, 135.0398, 135.2429, 135.7827, 136.3972, 137.1947, 138.0702, 138.6751, 139.3984, 140.0414, 140.7222, 141.3655, 141.7777, 142.3495, 143.3398, 144.6246, 145.7255, 146.9798, 147.8518, 148.4203, 149.1378, 149.7105, 150.2777, 150.7681, 151.3368, 152.0246, 152.5534, 153.3106, 154.1619, 155.1704, 157.1754, 158.8316, 160.3288, 161.8225, 163.417, 164.7778, 165.7041, 167.8735, 169.3755, 171.0168, 173.7187, 177.6018, 181.6882, 187.4093, 191.9621, 197.9857, 204.9622, 209.6414, 212.6967, 217.507, 223.3472, 230.0313, 235.5496, 239.4675, 243.4618, 246.6146, 249.734, 253.1245, 255.8553, 258.1288, 259.8069, 261.4982, 262.2751, 263.2001, 264.2001, 264.9347, 265.7699, 267.2728, 267.8286, 269.2026, 270.0261, 270.7131, 270.7926, 270.9941, 271.1283, 271.3225, 271.9303, 272.0029, 272.5711, 272.479, 272.5483, 272.8067, 273.0687, 273.0285, 273.4454, 273.3686, 273.4405, 273.2831, 272.6138, 272.9411, 103.0361, 102.2708, 101.8082, 101.6122, 101.5666, 101.5222, 101.4396, 101.432, 101.3845, 101.41, 101.7044, 103.9049, 107.3212, 109.6419, 110.618, 112.399, 114.6476, 115.966, 117.0682, 117.9726, 118.4546, 119.1334, 119.8885, 121.0288, 123.4719, 129.8989, 135.8431, 139.6448, 142.7624, 145.0349, 146.6238, 147.9886, 150.2946, 155.9004, 159.958, 162.5434, 164.7184, 169.3364, 178.3094, 185.4221, 190.8965, 197.0883, 212.2784, 226.9029, 241.5021, 250.7356, 256.102, 260.9407, 264.7889, 267.6385, 268.5046, 269.6416, 270.607, 271.2329, 272.0077, 272.4536, 272.7458, 273.5048, 273.2296, 273.2818, 96.8604, 96.4747, 96.6603, 96.6534, 96.7249, 96.8331, 97.1308, 97.1995, 97.4956, 98.2547, 98.8926, 99.4144, 99.7033, 99.7652, 99.8642, 100.1205, 101.2758, 102.4538, 104.9641, 107.5751, 109.2779, 110.7248, 112.0958, 113.4696, 114.9175, 115.9748, 118.053, 122.4135, 128.6701, 132.7799, 137.8979, 141.5471, 143.8999, 145.5656, 147.6261, 152.8154, 157.9403, 161.5384, 163.6583, 164.9434, 166.333, 168.4883, 173.3005, 178.69, 182.8189, 191.4581, 206.1119, 224.3167, 237.3205, 245.366, 252.0245, 258.0944, 263.5739, 266.4872, 268.7777, 269.9913, 270.7549, 271.8413, 272.448, 272.7374, 273.2827, 273.7304, 273.3509, 273.7351, 98.605, 97.7264, 97.3401, 97.1066, 97.0626, 97.1354, 97.1676, 97.3174, 97.6948, 98.3392, 98.7504, 99.0979, 100.2203, 102.5585, 104.2266, 105.5987, 107.2043, 108.6534, 110.8034, 112.4411, 113.5317, 114.4355, 115.9056, 118.1215, 119.635, 121.997, 125.3584, 128.2472, 131.4478, 135.0346, 138.4606, 141.1956, 143.4718, 144.9852, 148.0829, 153.825, 157.5161, 159.9736, 161.8098, 163.668, 167.8459, 173.3975, 177.3809, 186.9739, 203.3516, 217.1725, 229.6188, 237.1685, 242.2551, 246.4292, 250.4685, 258.2709, 264.0522, 267.7256, 269.6891, 271.2099, 272.2731, 273.3353, 274.2385, 274.3865, 274.5334, 274.7048, 88.6991, 89.2714, 89.6872, 89.8725, 90.1734, 90.7827, 91.1989, 91.1186, 91.1539, 91.6788, 92.2419, 92.9961, 93.9416, 94.9276, 95.3814, 95.4532, 95.9524, 96.3318, 96.6695, 97.0134, 97.2102, 97.754, 98.6068, 99.3693, 100.3609, 102.9875, 105.512, 107.3371, 108.7014, 109.534, 110.3662, 111.0463, 111.8934, 112.8796, 113.6348, 114.3876, 115.9214, 120.1416, 124.1191, 128.9309, 133.051, 136.131, 138.6397, 140.3412, 141.8162, 142.7181, 143.8503, 147.7885, 153.6134, 158.3733, 161.4628, 163.6563, 166.801, 171.6821, 176.3148, 183.8126, 196.1168, 208.3811, 216.4427, 225.3974, 232.4346, 239.052, 245.2603, 253.9012, 261.9194, 267.9997, 270.8156, 272.4863, 273.6227, 274.4424, 274.8847, 275.3942, 275.3052, 275.2478, 275.165, 275.0771, 275.2124, 78.5461, 77.8975, 77.8575, 77.9684, 78.1539, 78.301, 78.4108, 78.7514, 80.1238, 82.8778, 85.2483, 87.2699, 88.7917, 89.9287, 91.2189, 92.3961, 93.2617, 93.667, 94.0021, 94.4545, 95.4177, 96.2534, 96.5877, 96.2495, 95.8695, 95.7495, 95.9423, 96.1335, 96.477, 97.1636, 98.0328, 99.8483, 102.4996, 104.9758, 106.9202, 108.2524, 109.5959, 111.2403, 112.6864, 113.8252, 115.3546, 116.5694, 117.7007, 118.3772, 119.7485, 122.7547, 125.5643, 127.6897, 129.356, 131.1794, 133.6258, 137.1423, 140.4146, 145.7712, 151.8876, 156.8654, 158.9947, 161.1015, 163.683, 167.4813, 173.1871, 180.2405, 186.6733, 191.3736, 199.5234, 210.059, 223.8141, 237.0839, 244.8015, 250.5262, 256.3823, 261.2101, 264.4083, 266.5005, 267.287, 267.7322, 269.1219, 270.3822, 271.5348, 272.4581, 273.3163, 273.735, 273.9806, 274.1942, 82.7925, 82.4863, 82.9845, 83.862, 84.5422, 84.9968, 85.6835, 86.8682, 88.395, 89.5769, 90.2566, 90.9386, 91.5025, 91.9128, 92.3637, 92.814, 93.7368, 94.8506, 96.2288, 97.7509, 99.0131, 99.9237, 100.4922, 100.8636, 100.9678, 101.0338, 101.0618, 101.0904, 101.0879, 102.3997, 104.0461, 105.61, 107.1312, 107.8815, 108.328, 108.9006, 110.2156, 111.0438, 112.1496, 113.3636, 114.544, 115.9218, 117.7564, 119.4338, 121.9683, 124.4051, 126.386, 128.0585, 130.723, 136.2852, 145.49, 152.3542, 156.57, 158.6909, 159.8666, 160.413, 161.7226, 164.611, 166.7458, 169.9789, 174.2374, 179.0762, 185.8886, 191.6236, 197.4945, 203.8701, 209.5152, 214.0001, 225.0978, 236.5247, 245.9231, 252.8642, 257.2424, 261.7883, 264.8886, 266.4877, 267.7473, 268.5338, 268.9732, 269.6378, 269.8823, 270.5484, 271.3757, 271.3565, 88.3739, 88.3461, 88.9214, 89.2619, 89.686, 90.4127, 90.9412, 91.3541, 91.9995, 92.6838, 93.0959, 93.7849, 94.5447, 95.1458, 96.4457, 97.6649, 99.1945, 100.299, 101.0523, 101.6139, 102.1837, 102.6289, 102.8533, 103.1639, 103.8238, 104.2407, 104.4954, 104.5998, 104.8585, 105.3094, 105.6425, 107.1841, 108.5158, 109.3919, 110.0013, 110.4886, 110.7515, 111.1709, 111.3787, 111.9524, 112.6729, 113.3524, 114.1448, 115.2915, 117.5832, 118.7157, 121.0286, 123.6651, 125.2572, 126.3948, 127.3047, 127.981, 128.4291, 129.6851, 139.8878, 150.513, 156.2334, 159.8174, 160.4325, 161.1356, 163.9431, 167.1672, 172.495, 184.618, 194.6153, 202.3121, 207.6362, 212.2604, 216.9192, 221.1421, 223.9701, 230.9448, 239.9241, 245.8088, 251.3577, 257.0835, 260.8598, 263.895, 265.8571, 267.8158, 269.6341, 270.5574, 271.6326, 272.0374, 272.3588, 272.722, 272.6244, 59.9126, 60.7166, 62.6264, 63.9143, 65.2775, 65.989, 67.735, 69.0189, 70.7246, 72.7763, 74.0561, 75.3403, 76.6594, 77.9405, 79.2985, 80.386, 83.5577, 87.0195, 88.951, 90.7842, 92.755, 95.1218, 97.707, 98.913, 100.2813, 102.7843, 105.0007, 106.1372, 107.6547, 109.7754, 111.7921, 112.3212, 113.21, 114.88, 115.9894, 118.3562, 122.516, 126.1715, 128.0319, 131.0844, 149.6131, 161.6078, 167.3218, 176.3951, 194.7702, 212.2934, 222.9323, 227.6874, 227.5527, 234.6043, 246.2526, 256.194, 262.7636, 268.376, 271.2829, 272.6227, 273.0401, 273.0022, 56.9623, 56.8078, 57.7977, 58.7858, 59.8451, 60.75, 62.1139, 62.937, 63.149, 63.2853, 63.9572, 65.1641, 67.9876, 73.0973, 77.1248, 78.8588, 80.911, 82.7284, 86.1571, 89.1895, 90.6301, 91.5338, 92.2855, 93.0347, 94.2437, 95.993, 98.0496, 100.6285, 102.6151, 104.2369, 106.145, 107.8146, 109.8681, 111.9301, 113.7623, 115.2038, 116.1319, 118.2959, 123.6581, 128.4686, 131.4032, 140.01, 155.6012, 164.5, 170.1802, 179.716, 189.5214, 207.6327, 220.5697, 227.9658, 230.6632, 235.3312, 240.1127, 247.5982, 256.0879, 263.4666, 269.2109, 271.9763, 273.9438, 274.3612, 53.6852, 54.2559, 54.5536, 55.3177, 56.839, 57.3596, 57.6164, 58.18, 58.588, 59.2274, 59.9792, 61.4241, 62.5541, 63.9186, 66.1637, 68.1771, 72.024, 76.3743, 79.3439, 81.4221, 82.7863, 84.8396, 87.4209, 89.2732, 91.0892, 92.5595, 96.3295, 98.302, 97.7556, 96.3045, 97.4295, 98.7967, 100.4457, 102.3956, 104.867, 106.342, 109.1151, 111.429, 115.4545, 118.3402, 119.174, 119.4314, 120.6741, 123.8834, 126.8504, 128.6949, 130.5201, 132.8068, 140.8923, 148.5674, 157.1927, 170.0052, 181.5707, 194.2777, 204.7202, 211.4624, 220.8531, 231.837, 241.9405, 254.4899, 264.6883, 272.0302, 274.761, 275.4347, 275.584, 275.2763, 274.9223, 274.7921, 274.684, 49.2108, 49.0146, 48.9312, 48.8104, 48.54, 48.9548, 49.062, 49.6306, 50.2728, 51.413, 53.4309, 54.4884, 54.8583, 54.9624, 55.1809, 55.8953, 56.9158, 57.8202, 58.879, 61.702, 64.0916, 64.8395, 65.2887, 66.8836, 68.8587, 70.9074, 74.414, 77.0665, 78.8063, 81.616, 83.2028, 85.2529, 85.7849, 87.0755, 91.7133, 92.0847, 92.3796, 98.7642, 101.6576, 103.0301, 104.6212, 105.4418, 104.8928, 104.3433, 105.5959, 107.9855, 111.3073, 115.0809, 116.8991, 118.6675, 120.1482, 122.189, 124.0036, 125.8324, 129.0809, 132.3376, 135.4264, 139.7997, 149.7003, 163.8566, 174.3595, 182.6171, 192.0752, 197.6716, 200.7676, 208.9055, 218.2411, 226.0771, 233.6165, 242.0902, 251.6851, 260.1476, 267.1231, 269.5367, 270.4243, 271.0129, 271.4415, 271.7886, 272.4133, 272.8468, 40.8836, 40.6875, 40.5681, 40.4862, 40.4779, 40.3942, 40.4655, 41.2649, 42.7501, 43.4663, 44.1468, 44.8671, 46.2005, 46.956, 47.4464, 49.3101, 50.7109, 51.7713, 53.0998, 53.9673, 55.067, 56.2461, 58.1952, 60.0563, 62.1111, 63.706, 65.2997, 67.7711, 70.3946, 72.4838, 74.7207, 76.1196, 78.4394, 80.9497, 84.5653, 87.7521, 89.1074, 91.7988, 93.8417, 95.6309, 97.1864, 98.4259, 99.9424, 100.8456, 100.9612, 101.1919, 101.4165, 103.0649, 105.7951, 105.4183, 105.7023, 106.449, 108.73, 112.9224, 115.5389, 117.7522, 119.0846, 121.4068, 123.9126, 126.5366, 129.7946, 132.2741, 135.375, 137.8838, 139.9873, 143.8238, 152.1086, 155.7221, 158.3818, 162.5783, 167.7293, 172.8936, 180.2001, 189.8288, 206.2047, 225.9746, 231.7309, 236.1345, 240.997, 245.669, 250.6173, 260.9535, 265.6505, 268.8122, 271.1026, 271.8679, 41.1923, 41.3031, 42.1418, 43.286, 43.8495, 44.1854, 44.6762, 45.5502, 46.384, 46.9493, 47.5914, 48.0024, 48.3769, 49.0189, 50.0053, 51.3739, 52.7023, 53.6868, 54.4417, 55.12, 56.184, 57.281, 58.0, 59.841, 63.6543, 66.3517, 68.0947, 69.8783, 71.2007, 72.6017, 74.4255, 75.8228, 77.6058, 80.9139, 84.2933, 87.9045, 89.8054, 92.0846, 92.9907, 91.1265, 90.2741, 90.5636, 92.7701, 94.5111, 96.0374, 97.0982, 98.2435, 99.5581, 100.6283, 102.2997, 104.5825, 107.9302, 115.464, 121.5386, 125.2052, 127.1215, 127.2553, 126.4791, 125.2901, 126.472, 128.4101, 129.4558, 130.0503, 134.2048, 140.8144, 144.9724, 146.8733, 147.4612, 149.3221, 161.3065, 169.0868, 178.6013, 186.8777, 194.2755, 201.3965, 214.8778, 228.8367, 244.6635, 254.4287, 261.3243, 266.6216, 268.8421, 270.5023, 271.0456, 271.75, 272.0748, 272.3001, 27.7428, 27.8157, 28.386, 28.8401, 29.4877, 30.2067, 31.4237, 32.7216, 34.5133, 36.8808, 38.9045, 39.7341, 39.9503, 40.322, 41.96, 44.0564, 45.4596, 46.4839, 48.6903, 49.7467, 50.6141, 51.3624, 52.2655, 53.7786, 56.2125, 57.6485, 58.1667, 58.8469, 60.3672, 63.865, 65.9146, 70.4041, 75.3463, 78.5298, 87.8795, 88.4101, 88.5405, 90.6779, 93.3382, 95.4574, 96.8186, 98.0591, 99.1823, 101.9118, 104.0738, 106.256, 107.5099, 114.2405, 122.6885, 124.7446, 124.6421, 122.8354, 124.4634, 127.5645, 130.18, 131.6539, 133.3531, 135.1965, 139.8845, 150.2279, 158.4608, 173.3836, 193.8677, 212.0289, 225.3604, 234.2946, 241.6146, 254.6171, 268.8506, 272.8846, 274.2883, 274.9943}
    doxy_qc = 
      {1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1}
    time_gps = 
      {-999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0}
    longitude_gps = 
      {-999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0}
    latitude_gps = 
      {-999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0}
    gps_start_qc = 
      {0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0}
    gps_start_qc_tests = 
      {0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0}
    time_gps_end = 
      {1.6753619999999988E9, 1.6753650000000012E9, 1.6753680000000033E9, 1.6753709999999955E9, 1.6753741200000007E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754490000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754517000000033E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754544599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754571599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754598599999998E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.6754631600000043E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.675466639999998E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.6754699400000024E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.675473780000005E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754779199999995E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.6754821200000007E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.675486379999998E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754919000000012E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6754976599999998E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755039599999964E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.6755109800000005E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.675518360000003E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.6755259800000017E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9, 1.675534979999998E9}
    latitude_gps_end = 
      {38.3187, 38.3187, 38.3188, 38.3187, 38.3187, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2523, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2508, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2487, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2457, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2422, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2435, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2452, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2455, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2458, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.2468, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.247, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.248, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2497, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.2502, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.249, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.2478, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.245, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2655, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947, 38.2947}
    longitude_gps_end = 
      {-123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3467, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3543, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3623, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3693, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3762, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3832, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.3915, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4002, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4092, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.4182, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.428, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4382, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4555, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4742, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.4948, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5177, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5443, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5597, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762, -123.5762}
    gps_end_qc = 
      {0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0}
    gps_end_qc_tests = 
      {0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0}
    wmo_identifier =   "4801921"
    sensor_doxy = -127
    sensor_ctd = -127
    sensor_fchl = -127
    platform_model =   "Scripps Institution of Oceanography Spray glider"
    platform_serial_number =   "sp028"
    platform_meta = -127
    deployment_time = 
      {1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9, 1.675361294999998E9}
    deployment_latitude = 
      {38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187, 38.3187}
    deployment_longitude = 
      {-123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713, -123.0713}
}
